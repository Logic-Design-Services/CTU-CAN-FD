--------------------------------------------------------------------------------
-- 
-- CTU CAN FD IP Core 
-- Copyright (C) 2021-present Ondrej Ille
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to use, copy, modify, merge, publish, distribute the Component for
-- educational, research, evaluation, self-interest purposes. Using the
-- Component for commercial purposes is forbidden unless previously agreed with
-- Copyright holder.
-- 
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
-- 
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
-- 
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
-- 
-- -------------------------------------------------------------------------------
-- 
-- CTU CAN FD IP Core 
-- Copyright (C) 2015-2020 MIT License
-- 
-- Authors:
--     Ondrej Ille <ondrej.ille@gmail.com>
--     Martin Jerabek <martin.jerabek01@gmail.com>
-- 
-- Project advisors: 
-- 	Jiri Novak <jnovak@fel.cvut.cz>
-- 	Pavel Pisa <pisa@cmp.felk.cvut.cz>
-- 
-- Department of Measurement         (http://meas.fel.cvut.cz/)
-- Faculty of Electrical Engineering (http://www.fel.cvut.cz)
-- Czech Technical University        (http://www.cvut.cz/)
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to deal in the Component without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Component, and to permit persons to whom the
-- Component is furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
-- 
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
-- 
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
-- 
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- @TestInfoStart
--
-- @Purpose:
--  ERR_CAPT[ERR_POS] = ERC_POS_OVRL, Error code capture in Overload frame
--  feature test. 
--
-- @Verifies:
--  @1. Value of ERR_CAPT register when Error is detected inside Overload frame.
--
-- @Test sequence:
--  @1. Check that ERR_CAPT contains no error (post reset).
--  @2. Generate CAN frame and send it by DUT. Wait until intermission field
--      and force bus low (overload condition). Check that DUT transmitts
--      Overload frame. Wait for random number of bits (0-4) and force bus high
--      for one bit time. Check that DUT is transmitting Error frame. Read
--      Error code capture and check that error occured in Overload frame and
--      it was a bit error!
--
-- @TestInfoEnd
--------------------------------------------------------------------------------
-- Revision History:
--    12.01.2020   Created file
--------------------------------------------------------------------------------

Library ctu_can_fd_tb;
context ctu_can_fd_tb.ieee_context;
context ctu_can_fd_tb.rtl_context;
context ctu_can_fd_tb.tb_common_context;

use ctu_can_fd_tb.feature_test_agent_pkg.all;

package err_capt_ovr_frm_ftest is
    procedure err_capt_ovr_frm_ftest_exec(
        signal      chn             : inout  t_com_channel
    );
end package;


package body err_capt_ovr_frm_ftest is
    procedure err_capt_ovr_frm_ftest_exec(
        signal      chn             : inout  t_com_channel
    ) is
        -- Generated frames
        variable frame_1            :     t_ctu_frame;

        -- Node status
        variable stat_1             :     t_ctu_status;    

        variable wait_time          :     natural;
        variable frame_sent         :     boolean;
        variable err_capt           :     t_ctu_err_capt;
        variable mode_2             :     t_ctu_mode;
        
        variable pc_dbg             :     t_ctu_frame_field;
    begin

        -----------------------------------------------------------------------
        -- @1. Check that ERR_CAPT contains no error (post reset).
        -----------------------------------------------------------------------
        info_m("Step 1");
        
        ctu_get_err_capt(err_capt, DUT_NODE, chn);
        check_m(err_capt.err_pos = err_pos_other, "Reset of ERR_CAPT!");
        
        -----------------------------------------------------------------------
        -- @2. Generate CAN frame and send it by DUT. Wait until intermission
        --     field and force bus low (overload condition). Check that DUT
        --     transmitts Overload frame. Wait for random number of bits (0-4)
        --     and force bus high for one bit time. Check that DUT is
        --     transmitting Error frame. Read Error code capture and check that
        --     error occured in Overload frame and it was a bit error!
        -----------------------------------------------------------------------        
        generate_can_frame(frame_1);
        ctu_send_frame(frame_1, 1, DUT_NODE, chn, frame_sent);
        ctu_wait_frame_field(pc_deb_intermission, DUT_NODE, chn);
        wait for 20 ns;
        
        -- Cause overload condition
        force_bus_level(DOMINANT, chn);
        ctu_wait_sample_point(DUT_NODE, chn);
        wait for 20 ns; -- To be sure that opposite bit is sampled!
        release_bus_level(chn);
        
        ctu_get_curr_frame_field(pc_dbg, DUT_NODE, chn);
        check_m(pc_dbg = pc_deb_overload, "Overload frame transmitted!");
        
        rand_int_v(4, wait_time);
        info_m("Waiting for: " & integer'image(wait_time) & " bits!");
        for i in 1 to wait_time loop
            ctu_wait_sample_point(DUT_NODE, chn);
        end loop; 
        wait for 20 ns;

        -- Cause bit error in Overload frame!
        force_bus_level(RECESSIVE, chn);
        ctu_wait_sample_point(DUT_NODE, chn);
        wait for 20 ns; -- To be sure that opposite bit is sampled!
        release_bus_level(chn);

        ctu_get_status(stat_1, DUT_NODE, chn);
        check_m(stat_1.error_transmission, "Error frame is being transmitted!");

        ctu_get_err_capt(err_capt, DUT_NODE, chn);
        check_m(err_capt.err_type = can_err_bit, "Bit error detected!");
        check_m(err_capt.err_pos = err_pos_overload_frame,
                "Error detected in Overload frame!");
        
        -- For debug only to see waves properly!
        wait for 100 ns;

  end procedure;

end package body;
