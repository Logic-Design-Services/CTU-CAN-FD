--------------------------------------------------------------------------------
--
-- CTU CAN FD IP Core
-- Copyright (C) 2021-present Ondrej Ille
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to use, copy, modify, merge, publish, distribute the Component for
-- educational, research, evaluation, self-interest purposes. Using the
-- Component for commercial purposes is forbidden unless previously agreed with
-- Copyright holder.
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
--
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
--
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
--
-- -------------------------------------------------------------------------------
--
-- CTU CAN FD IP Core
-- Copyright (C) 2015-2020 MIT License
--
-- Authors:
--     Ondrej Ille <ondrej.ille@gmail.com>
--     Martin Jerabek <martin.jerabek01@gmail.com>
--
-- Project advisors:
-- 	Jiri Novak <jnovak@fel.cvut.cz>
-- 	Pavel Pisa <pisa@cmp.felk.cvut.cz>
--
-- Department of Measurement         (http://meas.fel.cvut.cz/)
-- Faculty of Electrical Engineering (http://www.fel.cvut.cz)
-- Czech Technical University        (http://www.cvut.cz/)
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to deal in the Component without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Component, and to permit persons to whom the
-- Component is furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
--
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
--
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
--
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- @TestInfoStart
--
-- @Purpose:
--  FDRF (Filter drop remote frame) feature test.
--
-- @Verifies:
--  @1. When SETTINGS[FDRF] is set, CTU CAN FD drops filters out RTR frames.
--  @1. When SETTINGS[FDRF] is NOT set, CTU CAN FD accepts RTR frames.
--
-- @Test sequence:
--  @1. Configure frame filters in DUT. Enable SETTINGS[FDRF]. Configure
--      filter A to accept any identifier (mask = all zeroes).4
--  @2. Send RTR frame by Test node. Wait until frame is sent and check that there
--      is no frame received by DUT.
--  @3. Disable SETTINGS[FDRF] in DUT.
--  @4. Send RTR frame by Test node. Wait until frame is sent and check that frame
--      is received by DUT.
--
-- @TestInfoEnd
--------------------------------------------------------------------------------
-- Revision History:
--    31.10.2020   Created file
--------------------------------------------------------------------------------

Library ctu_can_fd_tb;
context ctu_can_fd_tb.ieee_context;
context ctu_can_fd_tb.rtl_context;
context ctu_can_fd_tb.tb_common_context;

use ctu_can_fd_tb.feature_test_agent_pkg.all;

package mode_fdrf_ftest is
    procedure mode_fdrf_ftest_exec(
        signal      chn             : inout  t_com_channel
    );
end package;


package body mode_fdrf_ftest is
    procedure mode_fdrf_ftest_exec(
        signal      chn             : inout  t_com_channel
    ) is
        variable can_tx_frame       :       t_ctu_frame;
        variable can_rx_frame       :       t_ctu_frame;
        variable frame_sent         :       boolean := false;

        variable mode_1             :       t_ctu_mode := t_ctu_mode_rst_val;

        variable rx_buf_state       :       t_ctu_rx_buf_state;
        variable frames_equal       :       boolean := false;
        variable filt_A_cfg         :       t_ctu_mask_filt_cfg;
        variable filt_B_C_cfg       :       t_ctu_mask_filt_cfg;
        variable filter_range_cfg   :       t_ctu_ran_filt_cfg;

        variable hw_cfg             :       t_ctu_hw_cfg;
    begin

        ------------------------------------------------------------------------
        -- @1. Configure frame filters in DUT. Enable SETTINGS[FDRF].
        --     Configure filter A to accept any identifier (mask = all zeroes).
        ------------------------------------------------------------------------
        info_m("Step 1: Configure frame filters");

        -- Read HW config
        ctu_get_hw_config(hw_cfg, DUT_NODE, chn);

        if (hw_cfg.sup_filtA = false) then
            info_m("Skipping the test since sup_filtA=false");
            return;
        end if;

        mode_1.acceptance_filter := true;
        mode_1.fdrf := true;
        ctu_set_mode(mode_1, DUT_NODE, chn);

        -- Filter A (set mask to 0 - accept all frames)
        filt_A_cfg.ID_value := 0;
        filt_A_cfg.ID_mask := 0;
        filt_A_cfg.ident_type := BASE;
        filt_A_cfg.acc_CAN_2_0 := true;
        filt_A_cfg.acc_CAN_FD := true;
        ctu_set_mask_filter(filter_A, filt_A_cfg, DUT_NODE, chn);

        ------------------------------------------------------------------------
        -- @2. Send RTR frame by Test node. Wait until frame is sent and check
        --     that there is no frame received by DUT.
        ------------------------------------------------------------------------
        info_m("Step 2: Check that RTR frame is filtered when FDRF=1.");

        generate_can_frame(can_tx_frame);
        can_tx_frame.ident_type := BASE;
        can_tx_frame.frame_format := NORMAL_CAN;
        can_tx_frame.identifier := can_tx_frame.identifier mod 2048;
        can_tx_frame.rtr := RTR_FRAME;

        ctu_send_frame(can_tx_frame, 1, TEST_NODE, chn, frame_sent);
        ctu_wait_frame_sent(DUT_NODE, chn);

        ctu_get_rx_buf_state(rx_buf_state, DUT_NODE, chn);
        check_m(rx_buf_state.rx_frame_count = 0, "Frame filtered out!");

        ------------------------------------------------------------------------
        -- @3. Disable SETTINGS[FDRF] in DUT.
        ------------------------------------------------------------------------
        info_m("Step 3: Disable SETTINGS[FDRF]");

        mode_1.fdrf := false;
        ctu_set_mode(mode_1, DUT_NODE, chn);

        ------------------------------------------------------------------------
        -- @4. Send RTR frame by Test node. Wait until frame is sent and check
        --     that frame is received by DUT.
        ------------------------------------------------------------------------
        info_m("Step 4: Check that RTR frame is NOT filtered when FDRF=0.");

        generate_can_frame(can_tx_frame);
        can_tx_frame.ident_type := BASE;
        can_tx_frame.identifier := can_tx_frame.identifier mod 2048;
        can_tx_frame.rtr := RTR_FRAME;

        ctu_send_frame(can_tx_frame, 1, TEST_NODE, chn, frame_sent);
        ctu_wait_frame_sent(DUT_NODE, chn);

        ctu_get_rx_buf_state(rx_buf_state, DUT_NODE, chn);
        check_m(rx_buf_state.rx_frame_count = 1, "Frame NOT filtered out!");

  end procedure;

end package body;