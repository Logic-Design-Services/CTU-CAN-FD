--------------------------------------------------------------------------------
--
-- CTU CAN FD IP Core
-- Copyright (C) 2021-2023 Ondrej Ille
-- Copyright (C) 2023-     Logic Design Services Ltd.s
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to use, copy, modify, merge, publish, distribute the Component for
-- non-commercial purposes. Using the Component for commercial purposes is
-- forbidden unless previously agreed with Copyright holder.
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
--
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
--
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
--
-- -------------------------------------------------------------------------------
--
-- CTU CAN FD IP Core
-- Copyright (C) 2015-2020 MIT License
--
-- Authors:
--     Ondrej Ille <ondrej.ille@gmail.com>
--     Martin Jerabek <martin.jerabek01@gmail.com>
--
-- Project advisors:
-- 	Jiri Novak <jnovak@fel.cvut.cz>
-- 	Pavel Pisa <pisa@cmp.felk.cvut.cz>
--
-- Department of Measurement         (http://meas.fel.cvut.cz/)
-- Faculty of Electrical Engineering (http://www.fel.cvut.cz)
-- Czech Technical University        (http://www.cvut.cz/)
--
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to deal in the Component without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Component, and to permit persons to whom the
-- Component is furnished to do so, subject to the following conditions:
--
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
--
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
--
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
--
--------------------------------------------------------------------------------

library ctu_can_fd_tb;
context ctu_can_fd_tb.ieee_context;
use ctu_can_fd_tb.reference_test_agent_pkg.all;
use ctu_can_fd_tb.feature_test_agent_pkg.all;

package reference_data_set_5 is

constant C_reference_data_set_5 : t_reference_data_set := (
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 271377749,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 213586688,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 274361190,
         data => (x"66", x"24", x"a3", x"6a", x"0d", x"25", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 456290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 409293047,
         data => (x"02", x"5c", x"08", x"52", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1910 ns), ('0', 2010 ns), ('1', 465790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 147550791,
         data => (x"59", x"0c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 427290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1375,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1997,
         data => (x"af", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 451290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1382,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 289777569,
         data => (x"58", x"89", x"f2", x"b1", x"3a", x"54", x"9e", x"c8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 303290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 79
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1947,
         data => (x"d4", x"5e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1615,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 493310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 370972824,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  53542816,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 278211497,
         data => (x"78", x"68", x"39", x"c0", x"95", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 349290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 169178545,
         data => (x"c8", x"6c", x"f0", x"b3", x"09", x"17", x"cc", x"b5", x"05", x"23", x"1a", x"99", x"d5", x"1b", x"aa", x"89", x"3c", x"13", x"c7", x"50", x"2d", x"bf", x"b8", x"e5", x"00", x"4e", x"49", x"d1", x"b8", x"09", x"f7", x"82", x"75", x"e9", x"b5", x"fd", x"01", x"02", x"b4", x"85", x"26", x"4e", x"20", x"fb", x"69", x"4a", x"06", x"26", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 280790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 261
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1606,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 305888528,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 7990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 533670369,
         data => (x"b8", x"bf", x"ef", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 377310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1192,
         data => (x"18", x"3a", x"66", x"94", x"23", x"b0", x"9a", x"49", x"8e", x"e7", x"40", x"19", x"f4", x"70", x"0a", x"81", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 203310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 99
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 302152026,
         data => (x"36", x"5f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 423290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>  94152271,
         data => (x"41", x"64", x"7e", x"d8", x"1e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 373290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 293891906,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       108,
         data => (x"e3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 481290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>  42941565,
         data => (x"c4", x"4f", x"94", x"fb", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 461790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       572,
         data => (x"a9", x"be", x"b2", x"a7", x"97", x"d0", x"0d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 353290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1392,
         data => (x"c6", x"7c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 8110 ns), ('0', 1990 ns), ('1', 465290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>  78250076,
         data => (x"46", x"cb", x"56", x"8a", x"9a", x"ea", x"06", x"48", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 446310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 85
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1347,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 112801180,
         data => (x"d6", x"a2", x"24", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 411290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>  63066930,
         data => (x"a8", x"c5", x"8c", x"4a", x"11", x"52", x"95", x"67", x"dc", x"30", x"d2", x"e3", x"79", x"92", x"5b", x"3f", x"a1", x"fd", x"c4", x"e2", x"c7", x"e1", x"75", x"9e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 910 ns), ('0', 2010 ns), ('1', 382290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 147
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1788,
         data => (x"da", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 514810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>        95,
         data => (x"31", x"3d", x"62", x"18", x"99", x"93", x"6a", x"fc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 335290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 509402343,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 436307376,
         data => (x"f6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 409290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       934,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       644,
         data => (x"72", x"b8", x"03", x"af", x"1c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 417290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>  33823972,
         data => (x"3b", x"83", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 393310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 496304292,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1493,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 469290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 206950850,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 363591655,
         data => (x"3b", x"b1", x"50", x"d6", x"4d", x"19", x"85", x"d3", x"60", x"c0", x"57", x"80", x"47", x"7a", x"f7", x"de", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 2010 ns),
           ('1', 412790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 113
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 351365395,
         data => (x"66", x"e6", x"8d", x"8d", x"fc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 351310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier => 286888224,
         data => (x"3a", x"4b", x"2c", x"11", x"98", x"45", x"16", x"eb", x"26", x"d6", x"44", x"a6", x"1e", x"3e", x"1f", x"7d", x"dd", x"2d", x"65", x"98", x"8f", x"cb", x"00", x"1d", x"d8", x"fc", x"87", x"14", x"fb", x"20", x"ef", x"36", x"6b", x"9b", x"c6", x"84", x"60", x"dc", x"70", x"06", x"33", x"34", x"2d", x"52", x"72", x"4c", x"cf", x"50", x"79", x"b4", x"69", x"0a", x"00", x"69", x"a6", x"58", x"e5", x"2e", x"eb", x"e2", x"4f", x"5b", x"98", x"3a")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 212810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 311
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 495339026,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1738,
         data => (x"42", x"d7", x"57", x"91", x"a7", x"50", x"46", x"90", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 1990 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 488310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       668,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier => 515996068,
         data => (x"65", x"da", x"39", x"db", x"ba", x"f7", x"b2", x"77", x"a7", x"10", x"67", x"0d", x"1b", x"a9", x"64", x"f1", x"3b", x"8b", x"c2", x"01", x"1d", x"1c", x"c6", x"96", x"1d", x"e4", x"76", x"4d", x"ee", x"39", x"4b", x"54", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 990 ns), ('0', 990 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 351290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 183
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1761,
         data => (x"62", x"46", x"a4", x"73", x"ad", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 391290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       852,
         data => (x"91", x"a1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 465290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>  20076398,
         data => (x"54", x"fc", x"bd", x"cb", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 391310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 120909621,
         data => (x"99", x"99", x"30", x"69", x"96", x"93", x"af", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 319290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 290463189,
         data => (x"35", x"81", x"94", x"47", x"a2", x"57", x"d9", x"60", x"37", x"b3", x"b5", x"34", x"71", x"01", x"fd", x"9e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 165310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 117
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 265962876,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 304261753,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  70382612,
         data => (x"4c", x"6a", x"14", x"93", x"0e", x"ea", x"ec", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 450790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1114,
         data => (x"92", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      2015,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 495310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1178,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  98282528,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 478790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 376484906,
         data => (x"01", x"01", x"33", x"eb", x"ed", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 460810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 120473447,
         data => (x"a1", x"e9", x"38", x"d2", x"14", x"9e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 456790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  82897933,
         data => (x"84", x"c7", x"39", x"56", x"b6", x"da", x"11", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 319290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       284,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 168026287,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 451290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1494,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 520790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 118401948,
         data => (x"ac", x"88", x"a1", x"5b", x"0e", x"6a", x"94", x"64", x"a0", x"70", x"76", x"c3", x"b8", x"ad", x"67", x"82", x"18", x"f6", x"3a", x"25", x"95", x"01", x"77", x"18", x"e8", x"33", x"52", x"a3", x"82", x"aa", x"01", x"ae", x"33", x"23", x"0a", x"41", x"0d", x"9e", x"a6", x"ad", x"8e", x"9c", x"f0", x"c7", x"4a", x"58", x"4a", x"e1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns),
           ('1', 282290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 249
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       560,
         data => (x"7e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 449310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>  18561977,
         data => (x"b3", x"f7", x"12", x"e1", x"2c", x"b4", x"eb", x"6d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 301290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 81
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 302917872,
         data => (x"af", x"df", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 419310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1143,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 469310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 522211397,
         data => (x"e2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 474810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>  78948147,
         data => (x"c7", x"ad", x"46", x"a9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 397290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       752,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 336841113,
         data => (x"8c", x"9c", x"85", x"44", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 365310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       411,
         data => (x"b6", x"2d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 325202889,
         data => (x"04", x"04", x"00", x"4a", x"ad", x"d9", x"46", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 313290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>   8157127,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 451290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 262974930,
         data => (x"8b", x"01", x"04", x"ec", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 389290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1312,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       913,
         data => (x"7d", x"1a", x"73", x"48", x"48", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 389290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>        60,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier =>   4443965,
         data => (x"fc", x"cd", x"fc", x"7d", x"51", x"69", x"49", x"cd", x"9c", x"4c", x"f6", x"77", x"eb", x"70", x"8d", x"5f", x"6d", x"28", x"53", x"b5", x"70", x"a0", x"c3", x"fb", x"0f", x"d4", x"6d", x"79", x"16", x"7e", x"69", x"13", x"4c", x"66", x"90", x"1e", x"d0", x"59", x"eb", x"ec", x"25", x"62", x"e3", x"12", x"d2", x"72", x"f0", x"40", x"9a", x"c3", x"76", x"8a", x"64", x"b9", x"86", x"73", x"0f", x"74", x"6c", x"a4", x"f2", x"d6", x"37", x"40")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 212290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 319
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1345,
         data => (x"c9", x"fa", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  73775897,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 4110 ns), ('0', 2010 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  73687108,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier => 436098829,
         data => (x"e5", x"7d", x"f0", x"52", x"22", x"e3", x"a8", x"59", x"a3", x"66", x"a0", x"81", x"73", x"c0", x"ca", x"6e", x"07", x"76", x"4d", x"de", x"74", x"1e", x"28", x"b3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 375790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 147
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 153405743,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 416244385,
         data => (x"de", x"f5", x"d0", x"87", x"4f", x"f3", x"ed", x"6f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 299310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 79
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>       928,
         data => (x"b7", x"b7", x"9d", x"97", x"ab", x"3c", x"3f", x"5f", x"c5", x"f3", x"c7", x"44", x"1a", x"1e", x"c0", x"a6", x"72", x"2c", x"85", x"68", x"fc", x"8c", x"38", x"71", x"fa", x"a7", x"e6", x"5d", x"58", x"27", x"2d", x"11", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 383790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 169
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 326438002,
         data => (x"67", x"e9", x"cc", x"da", x"b1", x"11", x"f4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 343310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>       154,
         data => (x"a0", x"2b", x"fa", x"ad", x"e2", x"eb", x"a8", x"0b", x"d2", x"85", x"63", x"fa", x"32", x"74", x"d8", x"7d", x"9c", x"e3", x"84", x"83", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 435290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 125
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 290341281,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1963,
         data => (x"b1", x"10", x"be", x"2d", x"3d", x"21", x"19", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 387290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 119146503,
         data => (x"67", x"1d", x"84", x"40", x"1b", x"a1", x"a4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 315310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier =>         7,
         data => (x"f2", x"d2", x"57", x"44", x"06", x"c5", x"d6", x"b8", x"55", x"15", x"e5", x"92", x"37", x"7e", x"f7", x"63", x"6b", x"62", x"73", x"52", x"80", x"78", x"13", x"9b", x"1a", x"b7", x"ba", x"be", x"aa", x"2b", x"42", x"9d", x"fd", x"19", x"61", x"05", x"df", x"b8", x"3d", x"b4", x"cd", x"a2", x"c7", x"05", x"21", x"3f", x"e8", x"0d", x"a2", x"db", x"5f", x"23", x"54", x"f1", x"3e", x"6e", x"a9", x"f8", x"2e", x"d3", x"a4", x"ef", x"f1", x"22")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns), ('1', 470 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 1990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 250810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 323
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>       426,
         data => (x"e3", x"1e", x"5a", x"86", x"e5", x"de", x"28", x"26", x"c7", x"35", x"c8", x"a4", x"14", x"6b", x"f8", x"86", x"a9", x"e7", x"30", x"22", x"95", x"05", x"46", x"85", x"76", x"69", x"8f", x"49", x"10", x"f8", x"d5", x"f4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 2490 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 386810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 173
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 220791637,
         data => (x"a2", x"a3", x"d6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 910 ns), ('0', 2010 ns), ('1', 468790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       877,
         data => (x"f3", x"72", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 465290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1212,
         data => (x"27", x"e8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 465310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1130,
         data => (x"63", x"80", x"3d", x"d7", x"98", x"6d", x"52", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 385290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       172,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>  30153524,
         data => (x"42", x"ab", x"7d", x"9d", x"ce", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 373290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       294,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       747,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 372659619,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  33410409,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 2010 ns),
           ('1', 476790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>       241,
         data => (x"19", x"83", x"91", x"17", x"a1", x"df", x"b6", x"b0", x"56", x"40", x"b6", x"e9", x"1d", x"43", x"64", x"5c", x"51", x"9c", x"73", x"f6", x"c1", x"5d", x"33", x"62", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 2470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 418790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 133
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 392492404,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>  42554337,
         data => (x"75", x"3e", x"c0", x"2d", x"ee", x"96", x"6d", x"a5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9990 ns), ('0', 9990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 445810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 81
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 284296734,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1932,
         data => (x"b7", x"65", x"26", x"73", x"8e", x"7c", x"db", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 2010 ns), ('1', 357290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      2021,
         data => (x"0c", x"a9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 463290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1908,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1368,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 134870313,
         data => (x"5d", x"8d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 395290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1809,
         data => (x"2f", x"18", x"a6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 421290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1434,
         data => (x"83", x"e9", x"9b", x"da", x"ca", x"00", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 369310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 126806529,
         data => (x"2e", x"25", x"6d", x"f7", x"35", x"4a", x"85", x"7d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 6110 ns), ('0', 2010 ns), ('1', 295290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       904,
         data => (x"cf", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 481290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 492243113,
         data => (x"e1", x"e1", x"10", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 403310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 529560249,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>        24,
         data => (x"6e", x"5b", x"89", x"24", x"a5", x"8e", x"a1", x"b1", x"c7", x"d9", x"10", x"af", x"aa", x"13", x"5d", x"3d", x"71", x"83", x"20", x"53", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 432310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 125
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       444,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 469290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 196155477,
         data => (x"8f", x"a4", x"e5", x"98", x"c8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 351290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  43776534,
         data => (x"43", x"cc", x"9e", x"ed", x"e0", x"7b", x"ab", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 317290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       230,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 363340161,
         data => (x"1b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 441290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 255607595,
         data => (x"8b", x"2c", x"42", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 381310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>        13,
         data => (x"70", x"22", x"60", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 417290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       712,
         data => (x"d9", x"54", x"f9", x"eb", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 508970357,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1856,
         data => (x"1f", x"38", x"06", x"61", x"4f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>      1839,
         data => (x"c5", x"fb", x"db", x"48", x"58", x"e5", x"1d", x"b1", x"b9", x"17", x"9d", x"f7", x"c5", x"89", x"3a", x"15", x"11", x"00", x"3a", x"bd", x"5a", x"59", x"f5", x"60", x"ba", x"45", x"39", x"c8", x"68", x"d4", x"c6", x"2f", x"d1", x"a3", x"77", x"a9", x"09", x"15", x"da", x"c2", x"2c", x"79", x"3a", x"72", x"82", x"f3", x"87", x"93", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 321790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 241
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 240859830,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1177,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       953,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>  82495705,
         data => (x"af", x"13", x"54", x"5c", x"0c", x"0f", x"ce", x"0f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 297290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 442530817,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>       673,
         data => (x"08", x"c6", x"dc", x"27", x"bb", x"1a", x"8c", x"5f", x"a8", x"15", x"79", x"60", x"a6", x"2a", x"f2", x"fa", x"86", x"00", x"0a", x"55", x"8e", x"8d", x"aa", x"b0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1910 ns), ('0', 1990 ns),
           ('1', 418790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 145
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 390596686,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1657,
         data => (x"a4", x"e1", x"37", x"b0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 435290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 190400977,
         data => (x"6c", x"64", x"b3", x"e7", x"6a", x"33", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 361290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 402988910,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1753,
         data => (x"23", x"77", x"11", x"21", x"9d", x"2f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 403290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1045,
         data => (x"46", x"3c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 463310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 200001561,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 453310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 470622016,
         data => (x"2d", x"02", x"73", x"a0", x"86", x"20", x"b7", x"d6", x"c3", x"2f", x"e7", x"e4", x"4c", x"96", x"2a", x"4b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1910 ns), ('0', 1990 ns),
           ('1', 409810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 113
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 249922151,
         data => (x"04", x"49", x"07", x"62", x"03", x"18", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 10110 ns), ('0', 2010 ns),
           ('1', 357290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 141088054,
         data => (x"1b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 478790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 321414834,
         data => (x"f7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 2010 ns), ('1', 478290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1288,
         data => (x"77", x"9a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 510810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 453950928,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1650,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 275105525,
         data => (x"8b", x"0f", x"6d", x"b2", x"cb", x"8f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 456790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1898,
         data => (x"e7", x"f4", x"d1", x"60", x"8f", x"0c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 371290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 149825860,
         data => (x"99", x"8e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 425290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 486277984,
         data => (x"84", x"0f", x"28", x"94", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 361310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 476476923,
         data => (x"a0", x"14", x"59", x"03", x"fc", x"4f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 329290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 499730402,
         data => (x"2a", x"32", x"3e", x"8f", x"cb", x"4c", x"94", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 315290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 354226560,
         data => (x"61", x"d4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 395310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 196640711,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier => 218555842,
         data => (x"fb", x"ac", x"51", x"d8", x"0b", x"32", x"8a", x"b5", x"64", x"c8", x"45", x"30", x"95", x"59", x"c0", x"f3", x"aa", x"ed", x"57", x"0c", x"42", x"4f", x"6a", x"71", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 378790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 157
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  62697668,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 211055161,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>      1388,
         data => (x"04", x"7d", x"83", x"b4", x"13", x"dc", x"f4", x"87", x"88", x"63", x"5e", x"14", x"a5", x"ae", x"7f", x"18", x"56", x"d4", x"0d", x"75", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 490 ns), ('1', 910 ns), ('0', 2010 ns), ('1', 435290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 127
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>  51491510,
         data => (x"fd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 364048238,
         data => (x"22", x"d8", x"a9", x"56", x"ec", x"87", x"4b", x"f3", x"8f", x"ae", x"52", x"a3", x"55", x"80", x"a2", x"6d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 171310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 121
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 159233955,
         data => (x"59", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 441290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  48261017,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1383,
         data => (x"79", x"ed", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 512810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 440584786,
         data => (x"04", x"6d", x"ab", x"27", x"c2", x"ac", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 355290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       413,
         data => (x"cf", x"e4", x"82", x"2e", x"83", x"b8", x"0b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 349290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 151430628,
         data => (x"21", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 411290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 362596385,
         data => (x"d0", x"20", x"7f", x"3e", x"4b", x"a6", x"80", x"f7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 291310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       603,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       740,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       614,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1457,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 189425717,
         data => (x"85", x"cd", x"5f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 405310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 529523340,
         data => (x"52", x"52", x"d6", x"9e", x"6c", x"32", x"98", x"89", x"c5", x"1d", x"ee", x"2f", x"a6", x"3b", x"b2", x"51", x"e8", x"bc", x"0f", x"db", x"c2", x"9d", x"ef", x"c7", x"ea", x"ce", x"74", x"b9", x"a5", x"92", x"b7", x"f8", x"64", x"0e", x"97", x"51", x"40", x"af", x"da", x"86", x"cc", x"c9", x"b5", x"73", x"85", x"e8", x"44", x"ed", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 510 ns), ('1', 970 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1410 ns), ('0', 2010 ns), ('1', 279790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 259
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>       632,
         data => (x"39", x"b0", x"db", x"08", x"25", x"15", x"ae", x"37", x"4c", x"27", x"9c", x"d9", x"3e", x"ed", x"1b", x"ed", x"48", x"21", x"3a", x"13", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 434290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 115
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 125943433,
         data => (x"06", x"65", x"c3", x"4f", x"4e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 373310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1908,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  15169073,
         data => (x"66", x"78", x"4a", x"a4", x"66", x"e4", x"12", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 450310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>      1878,
         data => (x"78", x"5a", x"1c", x"69", x"df", x"81", x"2d", x"2f", x"cf", x"61", x"b8", x"4e", x"ef", x"ca", x"73", x"94", x"8a", x"50", x"04", x"71", x"c8", x"4e", x"16", x"af", x"33", x"a8", x"5f", x"39", x"74", x"21", x"16", x"ed", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1910 ns), ('0', 1990 ns),
           ('1', 387310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 177
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       934,
         data => (x"84", x"0a", x"82", x"e5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 429310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 458859627,
         data => (x"e9", x"97", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 2010 ns), ('1', 474790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       703,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       676,
         data => (x"2a", x"bc", x"0d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 449290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier => 411549028,
         data => (x"e2", x"a4", x"86", x"6d", x"a6", x"eb", x"30", x"f7", x"41", x"bd", x"3c", x"2c", x"55", x"d0", x"9a", x"5f", x"ad", x"d7", x"fe", x"3b", x"c8", x"47", x"27", x"f3", x"83", x"b4", x"b3", x"2e", x"bc", x"26", x"30", x"20", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 346790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 175
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 169905386,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 482790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1139,
         data => (x"8e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 483290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1711,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 4110 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 312310027,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1560,
         data => (x"a6", x"f7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 435290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>        31,
         data => (x"a4", x"d2", x"2e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 447310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 252894402,
         data => (x"20", x"ac", x"d6", x"c8", x"da", x"fa", x"c9", x"09", x"59", x"14", x"fc", x"df", x"d0", x"75", x"1b", x"42", x"1c", x"93", x"59", x"72", x"2b", x"3b", x"fe", x"50", x"8d", x"ac", x"b1", x"4a", x"3e", x"8e", x"2b", x"dd", x"ba", x"82", x"26", x"95", x"fc", x"70", x"1e", x"56", x"84", x"1c", x"37", x"55", x"91", x"d1", x"18", x"2e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 282310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 255
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1287,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       411,
         data => (x"84", x"8a", x"21", x"2f", x"68", x"db", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 375310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>  89729591,
         data => (x"10", x"85", x"04", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 381290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1538,
         data => (x"f0", x"eb", x"f3", x"62", x"0c", x"84", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 369310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 522594252,
         data => (x"77", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 437290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 210164319,
         data => (x"f4", x"ad", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 425290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1334,
         data => (x"e1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 481310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1793,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1276,
         data => (x"d9", x"23", x"3a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 2010 ns),
           ('1', 447290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 248891220,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 7990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1375,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       920,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1323,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 520790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 290710656,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 269069533,
         data => (x"f0", x"a0", x"4c", x"f3", x"1f", x"4c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 331310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 336899866,
         data => (x"f3", x"8a", x"fd", x"69", x"e0", x"e5", x"57", x"19", x"4d", x"69", x"6e", x"0e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 231290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 95
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 212852086,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 301125443,
         data => (x"21", x"33", x"f5", x"6d", x"76", x"19", x"d2", x"07", x"2b", x"46", x"11", x"a9", x"b0", x"f1", x"8f", x"87", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 167290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 109
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1465,
         data => (x"4c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1778,
         data => (x"20", x"cd", x"90", x"77", x"ee", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 385290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 281633672,
         data => (x"2e", x"41", x"b1", x"f4", x"53", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 373310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 409920991,
         data => (x"50", x"47", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 470290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       744,
         data => (x"36", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 483290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 324120517,
         data => (x"18", x"e9", x"69", x"5b", x"d7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 351290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1077,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       305,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1707,
         data => (x"57", x"0a", x"4f", x"c1", x"3c", x"05", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 399290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 407012324,
         data => (x"a3", x"f1", x"4c", x"7f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 387290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 255039147,
         data => (x"6c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 441310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 193333472,
         data => (x"08", x"f5", x"35", x"c7", x"12", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 349290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 362206604,
         data => (x"e5", x"63", x"f5", x"72", x"6b", x"d8", x"95", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 343290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 518578541,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 459310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       683,
         data => (x"a8", x"2f", x"26", x"23", x"b6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 417310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 208535021,
         data => (x"50", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 2010 ns), ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1629,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>  95438337,
         data => (x"de", x"52", x"13", x"06", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 393310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 498969708,
         data => (x"59", x"ec", x"03", x"00", x"10", x"39", x"1b", x"e8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 2010 ns),
           ('1', 446290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       373,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 495310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 391506499,
         data => (x"b5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 443310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 312889362,
         data => (x"45", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 476790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier =>      1161,
         data => (x"57", x"2c", x"f3", x"d9", x"ab", x"84", x"14", x"c6", x"6d", x"4c", x"90", x"3b", x"d4", x"69", x"3c", x"3b", x"37", x"d4", x"f5", x"6c", x"ee", x"de", x"1f", x"e6", x"99", x"e4", x"65", x"dc", x"67", x"b7", x"65", x"3e", x"63", x"d8", x"98", x"0f", x"dc", x"ac", x"56", x"c9", x"f8", x"e6", x"05", x"4d", x"cf", x"42", x"08", x"07", x"96", x"7d", x"73", x"85", x"5c", x"12", x"ec", x"f5", x"f6", x"52", x"53", x"de", x"89", x"b8", x"9c", x"ed")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 255290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 309
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1168,
         data => (x"52", x"b8", x"5a", x"39", x"3e", x"27", x"09", x"80", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 337290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>       943,
         data => (x"9c", x"89", x"16", x"89", x"00", x"8c", x"db", x"53", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 341310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 432732787,
         data => (x"1c", x"bd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 425290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1945,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 469290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 370419156,
         data => (x"02", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 439290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 506946207,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1990,
         data => (x"9a", x"99", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 510790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       386,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       474,
         data => (x"ec", x"43", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 465310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 386134970,
         data => (x"03", x"55", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 393310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1454,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       956,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       136,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       297,
         data => (x"ed", x"ba", x"64", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 419290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 255774785,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 8090 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 255695300,
         data => (x"22", x"09", x"3a", x"45", x"e9", x"b6", x"a7", x"53", x"4e", x"23", x"17", x"6b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 432310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 99
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       162,
         data => (x"8e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>  42169467,
         data => (x"be", x"d8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 470290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1109,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 498169324,
         data => (x"36", x"e6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 399290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>  21175328,
         data => (x"20", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 437290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 379164171,
         data => (x"45", x"5b", x"fa", x"b7", x"e3", x"30", x"f6", x"3d", x"45", x"0b", x"e8", x"8e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 233290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 97
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 392181250,
         data => (x"ab", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       449,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 8110 ns), ('0', 1990 ns),
           ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 17
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1692,
         data => (x"03", x"99", x"2f", x"c7", x"74", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 415310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1128,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>       779,
         data => (x"cf", x"5e", x"29", x"e9", x"ed", x"54", x"ba", x"64", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 343290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       648,
         data => (x"5d", x"6d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 435290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1842,
         data => (x"7c", x"47", x"a8", x"55", x"23", x"9f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 373290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>        61,
         data => (x"f0", x"48", x"9c", x"db", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       991,
         data => (x"2b", x"aa", x"1f", x"ba", x"08", x"8d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 397290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>      1275,
         data => (x"91", x"8c", x"39", x"67", x"2f", x"d8", x"d2", x"f2", x"f9", x"bd", x"e4", x"ea", x"06", x"81", x"46", x"3c", x"72", x"dc", x"d6", x"3b", x"08", x"81", x"5a", x"42", x"0a", x"67", x"e9", x"72", x"7c", x"2e", x"83", x"8e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 383310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 169
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1824,
         data => (x"48", x"5c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 510790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 105785360,
         data => (x"43", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 437290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 302736382,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 392751963,
         data => (x"2b", x"32", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 399290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 500202263,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 482790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 480727501,
         data => (x"f1", x"7b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 397290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>       423,
         data => (x"8e", x"84", x"3c", x"57", x"ba", x"59", x"f6", x"aa", x"fd", x"97", x"75", x"64", x"43", x"a8", x"35", x"60", x"d7", x"33", x"02", x"15", x"ec", x"de", x"c7", x"90", x"51", x"c2", x"10", x"52", x"c4", x"d1", x"4d", x"53", x"56", x"09", x"2a", x"90", x"62", x"a0", x"3c", x"df", x"39", x"b1", x"44", x"fb", x"d9", x"f8", x"5c", x"b1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 319790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 245
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 203650966,
         data => (x"0e", x"2a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 421290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1104,
         data => (x"8b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 451290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>        38,
         data => (x"f2", x"1b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 510810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier => 376138707,
         data => (x"bf", x"e9", x"ba", x"38", x"46", x"ec", x"e4", x"a4", x"b2", x"7f", x"e1", x"41", x"29", x"70", x"92", x"e3", x"d0", x"28", x"6f", x"7f", x"12", x"51", x"b8", x"a6", x"45", x"53", x"5b", x"73", x"cd", x"49", x"54", x"0d", x"b2", x"8f", x"46", x"78", x"7c", x"aa", x"1d", x"ae", x"2a", x"fe", x"ef", x"d3", x"ee", x"82", x"b7", x"c0", x"ab", x"a6", x"40", x"3d", x"f8", x"78", x"63", x"bd", x"cb", x"be", x"31", x"1a", x"08", x"86", x"a6", x"3a")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 214310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 321
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 387072397,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 432614657,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 116942713,
         data => (x"de", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 342243717,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 169900567,
         data => (x"9f", x"c7", x"e1", x"c5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 391290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>  63005345,
         data => (x"ca", x"07", x"4a", x"8c", x"57", x"fa", x"23", x"97", x"2e", x"ef", x"97", x"0e", x"64", x"58", x"2b", x"51", x"92", x"2b", x"fb", x"18", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 510 ns), ('1', 970 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 2010 ns), ('1', 397790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 135
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 463057076,
         data => (x"fc", x"36", x"b2", x"af", x"6c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 8110 ns), ('0', 1990 ns),
           ('1', 375310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>  30992421,
         data => (x"cb", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 474790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       512,
         data => (x"fa", x"3d", x"7f", x"54", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 429310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 230355219,
         data => (x"7e", x"fe", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 423290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 157394943,
         data => (x"68", x"91", x"e2", x"d4", x"4d", x"5d", x"c7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1390 ns), ('0', 2010 ns), ('1', 450790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1897,
         data => (x"76", x"02", x"ab", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1390 ns), ('0', 2010 ns), ('1', 508290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 280262697,
         data => (x"fa", x"2c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 9990 ns),
           ('1', 8110 ns), ('0', 2010 ns), ('1', 419290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>  97737560,
         data => (x"df", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 478810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1981,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       761,
         data => (x"7e", x"b7", x"82", x"51", x"48", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 385290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1897,
         data => (x"1e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 133759789,
         data => (x"e1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 8110 ns), ('0', 1990 ns), ('1', 437290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1635,
         data => (x"9a", x"79", x"67", x"79", x"ee", x"0e", x"24", x"41", x"fc", x"a2", x"78", x"80", x"f3", x"c0", x"f9", x"c6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 203310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 91
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 250836064,
         data => (x"90", x"eb", x"74", x"82", x"cd", x"7c", x"ac", x"9b", x"e3", x"c0", x"37", x"dc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 430290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 91
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1111,
         data => (x"0c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       626,
         data => (x"46", x"2d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 512790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 226644013,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 171230777,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 459310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 295121442,
         data => (x"8b", x"d9", x"da", x"b3", x"89", x"a5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 456790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>       546,
         data => (x"38", x"51", x"c0", x"fd", x"fd", x"f2", x"f8", x"91", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 910 ns), ('0', 2010 ns), ('1', 485790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1891,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier => 266075672,
         data => (x"a9", x"70", x"0e", x"03", x"ca", x"c1", x"8c", x"70", x"ab", x"e9", x"23", x"c8", x"bf", x"da", x"99", x"00", x"d9", x"18", x"f2", x"d2", x"a9", x"ef", x"99", x"e3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 990 ns), ('1', 990 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 374790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 141
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>      1644,
         data => (x"af", x"44", x"4b", x"9f", x"52", x"4e", x"6a", x"14", x"5a", x"da", x"bf", x"44", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 471790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 95
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 188680909,
         data => (x"03", x"33", x"3a", x"75", x"86", x"e3", x"66", x"20", x"47", x"70", x"3a", x"84", x"b1", x"db", x"34", x"f5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 169310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 111
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 443382778,
         data => (x"5c", x"ce", x"98", x"1c", x"93", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 349290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 342477661,
         data => (x"9a", x"24", x"01", x"10", x"aa", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 377290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 329810504,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 204406697,
         data => (x"0f", x"88", x"b7", x"58", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 361310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>        15,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 493290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1266,
         data => (x"96", x"3c", x"91", x"3b", x"bc", x"21", x"65", x"21", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 343290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>  74821517,
         data => (x"fc", x"97", x"98", x"e0", x"a7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 347310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       106,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1575,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 9990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 8110 ns), ('0', 1990 ns),
           ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 17
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>        37,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 117856501,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>      1868,
         data => (x"e2", x"5d", x"23", x"fa", x"3e", x"ca", x"9c", x"57", x"4a", x"ba", x"67", x"fd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 273310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 89
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 354073724,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 120332402,
         data => (x"b8", x"a5", x"f9", x"34", x"b9", x"06", x"e0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 333290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       597,
         data => (x"3f", x"35", x"fd", x"db", x"8d", x"c7", x"16", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns),
           ('1', 491790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 429026608,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 429310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 231262438,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>        19,
         data => (x"53", x"59", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 435290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       419,
         data => (x"e9", x"2b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 328195180,
         data => (x"f1", x"28", x"20", x"38", x"e4", x"1a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 353310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 388515565,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier => 358992794,
         data => (x"3b", x"b2", x"3a", x"22", x"e5", x"2d", x"99", x"dd", x"96", x"c4", x"13", x"b6", x"ee", x"25", x"62", x"61", x"cc", x"83", x"99", x"b1", x"1d", x"9b", x"44", x"f8", x"e3", x"b7", x"3a", x"a4", x"92", x"99", x"86", x"4e", x"cc", x"c0", x"ef", x"32", x"6e", x"89", x"10", x"05", x"4e", x"a3", x"3b", x"3e", x"48", x"1e", x"9f", x"15", x"a1", x"b8", x"46", x"3e", x"54", x"0a", x"b6", x"b7", x"c1", x"f0", x"5d", x"d4", x"0a", x"63", x"a2", x"56")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 216790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 323
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1963,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 469290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1663,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>      1639,
         data => (x"12", x"80", x"de", x"cf", x"54", x"e8", x"86", x"8c", x"ab", x"77", x"69", x"80", x"02", x"cc", x"23", x"d7", x"70", x"35", x"61", x"03", x"51", x"fa", x"9a", x"3b", x"37", x"6d", x"e3", x"bc", x"de", x"2b", x"d5", x"70", x"2b", x"b5", x"41", x"80", x"9e", x"c7", x"0d", x"c9", x"bf", x"76", x"c9", x"41", x"43", x"6c", x"19", x"33", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 490 ns),
           ('1', 910 ns), ('0', 2010 ns), ('1', 320290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 243
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 319577369,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>       694,
         data => (x"69", x"1d", x"3d", x"bf", x"8d", x"69", x"f4", x"4e", x"e9", x"13", x"96", x"76", x"dd", x"d5", x"ec", x"27", x"17", x"af", x"94", x"af", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 2010 ns), ('1', 436790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 125
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 480326201,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       134,
         data => (x"e9", x"36", x"c5", x"27", x"f5", x"54", x"10", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 353290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 177001262,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       925,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 142619188,
         data => (x"cd", x"7f", x"88", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 407290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       295,
         data => (x"9c", x"38", x"a2", x"62", x"de", x"99", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 375290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       644,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 469310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 470754481,
         data => (x"b5", x"e0", x"c5", x"42", x"77", x"1b", x"31", x"45", x"1b", x"b9", x"bb", x"ba", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 2010 ns),
           ('1', 430290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 97
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1572,
         data => (x"c9", x"2b", x"a0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 449290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 238918451,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 248873281,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 478790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       324,
         data => (x"9e", x"4f", x"fb", x"64", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 2010 ns), ('1', 405290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>       951,
         data => (x"2a", x"4b", x"2a", x"6b", x"15", x"55", x"0c", x"78", x"36", x"9b", x"5f", x"71", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 275290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 91
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      2007,
         data => (x"ab", x"70", x"b5", x"de", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>  76690319,
         data => (x"18", x"eb", x"59", x"bc", x"cd", x"83", x"87", x"f7", x"6f", x"1d", x"cc", x"fa", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 235290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 83
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 492097139,
         data => (x"ac", x"3c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 427310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 448596292,
         data => (x"81", x"3c", x"40", x"56", x"6a", x"77", x"8f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 339290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 200140018,
         data => (x"ec", x"c7", x"a8", x"db", x"e4", x"75", x"57", x"f9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 510 ns), ('1', 970 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1410 ns), ('0', 2010 ns), ('1', 447790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1017,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>      1200,
         data => (x"b4", x"78", x"b7", x"75", x"4e", x"a2", x"ec", x"de", x"a5", x"cf", x"48", x"64", x"81", x"b4", x"2c", x"2a", x"91", x"90", x"20", x"e8", x"8a", x"19", x"57", x"f8", x"05", x"72", x"24", x"a3", x"a1", x"1a", x"9f", x"d6", x"12", x"d6", x"4c", x"61", x"79", x"b8", x"40", x"9e", x"88", x"08", x"04", x"0a", x"bc", x"af", x"b4", x"cd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 318810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 253
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1411,
         data => (x"0d", x"45", x"f1", x"7f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1977,
         data => (x"f8", x"16", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 433310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier => 484559125,
         data => (x"37", x"25", x"05", x"3f", x"29", x"8f", x"7b", x"59", x"44", x"c9", x"9a", x"98", x"00", x"e5", x"85", x"0e", x"2b", x"77", x"0d", x"14", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 398290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 139
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 131660619,
         data => (x"ad", x"d0", x"eb", x"a4", x"d7", x"68", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 454810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1646,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 520790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1326,
         data => (x"1a", x"5a", x"df", x"00", x"5f", x"6d", x"ab", x"d6", x"7a", x"3f", x"65", x"2a", x"d6", x"a8", x"51", x"04", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 203290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 113
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 275004150,
         data => (x"04", x"4e", x"14", x"9d", x"f3", x"91", x"34", x"73", x"d2", x"13", x"8d", x"ac", x"f2", x"0d", x"0c", x"df", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 7990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 415310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 101
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       215,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       611,
         data => (x"6b", x"13", x"fc", x"bb", x"b9", x"81", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 399290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1915,
         data => (x"d2", x"f0", x"32", x"e6", x"fd", x"df", x"59", x"0c", x"eb", x"3a", x"44", x"4f", x"15", x"bc", x"97", x"99", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1990 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 103
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       258,
         data => (x"83", x"dd", x"30", x"3d", x"de", x"ba", x"8a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 375310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>  68329650,
         data => (x"1d", x"b7", x"27", x"fc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 361290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 102809521,
         data => (x"38", x"df", x"34", x"cf", x"79", x"c0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 455790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 312947550,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 145772879,
         data => (x"33", x"5d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 427310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1765,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>         0,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 465310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1807,
         data => (x"22", x"27", x"1b", x"e2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 504310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>  90306990,
         data => (x"85", x"cd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 421290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 434584517,
         data => (x"79", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1690 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 476810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>  45398820,
         data => (x"56", x"58", x"ce", x"cc", x"f6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 375290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 280722419,
         data => (x"f5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 476290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1380,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>      1638,
         data => (x"ad", x"1b", x"a5", x"6f", x"94", x"0d", x"60", x"a8", x"2f", x"b7", x"fe", x"88", x"86", x"4b", x"fe", x"97", x"85", x"4e", x"4b", x"e0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 127
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 271931821,
         data => (x"e3", x"80", x"ae", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81900 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 467810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       227,
         data => (x"2e", x"4b", x"c4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 449290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       784,
         data => (x"6d", x"73", x"e9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 447290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier => 488633551,
         data => (x"4d", x"9f", x"05", x"67", x"3f", x"3f", x"53", x"a3", x"bf", x"03", x"d0", x"d4", x"8b", x"2c", x"05", x"3a", x"f7", x"c9", x"76", x"24", x"b7", x"61", x"87", x"a4", x"55", x"71", x"dc", x"48", x"72", x"9b", x"09", x"3f", x"3b", x"8d", x"26", x"f9", x"cc", x"7a", x"9d", x"0c", x"fc", x"ee", x"e0", x"08", x"1b", x"65", x"42", x"92", x"30", x"38", x"b6", x"67", x"1a", x"bd", x"0c", x"ee", x"2f", x"e8", x"37", x"22", x"84", x"bf", x"e0", x"3f")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 2490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1910 ns), ('0', 1990 ns), ('1', 210810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 315
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier => 114431156,
         data => (x"57", x"a5", x"7e", x"c5", x"07", x"06", x"61", x"6c", x"49", x"f3", x"1c", x"01", x"ab", x"83", x"9a", x"e8", x"8f", x"89", x"98", x"79", x"40", x"ba", x"7d", x"00", x"1b", x"3d", x"cc", x"a2", x"f6", x"66", x"a4", x"cd", x"0d", x"a2", x"94", x"14", x"a9", x"f5", x"80", x"72", x"69", x"9d", x"f2", x"94", x"21", x"8e", x"7e", x"31", x"97", x"17", x"2a", x"d8", x"51", x"27", x"58", x"6c", x"64", x"26", x"10", x"5b", x"0c", x"34", x"2a", x"19")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1970 ns), ('0', 2510 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 990 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 215810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 313
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>        21,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1049,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 115093131,
         data => (x"8c", x"c7", x"c6", x"e4", x"19", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 371290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 478108268,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 136048549,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 3990 ns), ('1', 4110 ns), ('0', 2010 ns), ('1', 451290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>       713,
         data => (x"4a", x"e3", x"93", x"67", x"ae", x"f8", x"1a", x"1a", x"6d", x"ca", x"b7", x"79", x"92", x"7e", x"dd", x"2b", x"ec", x"9a", x"b0", x"41", x"fd", x"c4", x"ef", x"ec", x"0e", x"c8", x"f4", x"2e", x"5f", x"aa", x"ce", x"a9", x"0e", x"e1", x"11", x"bc", x"5b", x"ab", x"57", x"48", x"f5", x"0f", x"41", x"09", x"0d", x"1f", x"b3", x"fa", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 319790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 249
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1216,
         data => (x"ab", x"a3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 435310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 198417113,
         data => (x"44", x"b4", x"fc", x"53", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 464290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1418,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 331525782,
         data => (x"38", x"83", x"1a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 381310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>      1675,
         data => (x"0b", x"7a", x"65", x"ae", x"b1", x"59", x"c7", x"97", x"ac", x"0d", x"4d", x"29", x"df", x"64", x"b6", x"6f", x"d5", x"ef", x"d6", x"10", x"1f", x"4c", x"0b", x"57", x"4f", x"a4", x"c2", x"4d", x"f7", x"13", x"07", x"82", x"0d", x"eb", x"b1", x"bf", x"c4", x"79", x"57", x"f0", x"06", x"24", x"1a", x"65", x"08", x"51", x"d5", x"dd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 2490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 317310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 241
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1189,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1367,
         data => (x"16", x"15", x"0e", x"9d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  33304301,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 451310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 526105968,
         data => (x"56", x"5a", x"2f", x"de", x"2b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 371310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       646,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1107,
         data => (x"40", x"fc", x"88", x"55", x"8a", x"26", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 2010 ns), ('1', 371290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>        32,
         data => (x"7d", x"79", x"32", x"bd", x"42", x"89", x"18", x"f0", x"68", x"43", x"75", x"a4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 271290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 85
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 429740933,
         data => (x"f2", x"7e", x"41", x"33", x"fa", x"49", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 329290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  48126226,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 444189509,
         data => (x"df", x"d9", x"67", x"e8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 391310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>        44,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 263059624,
         data => (x"43", x"38", x"dc", x"05", x"6b", x"d8", x"4e", x"f3", x"de", x"3e", x"e8", x"0b", x"dc", x"15", x"b7", x"f8", x"b9", x"17", x"d3", x"21", x"00", x"c4", x"f9", x"50", x"7a", x"c7", x"c6", x"5d", x"bb", x"0c", x"bc", x"7f", x"44", x"19", x"84", x"2f", x"71", x"d2", x"a2", x"50", x"11", x"8b", x"5b", x"ed", x"20", x"93", x"67", x"5a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 276290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 237
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1312,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1376,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 8090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>        15,
         data => (x"91", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 481290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 274357989,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 480790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 199946022,
         data => (x"4e", x"0f", x"5f", x"b5", x"e8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1910 ns), ('0', 1990 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>        65,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 17
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 148542395,
         data => (x"42", x"8e", x"c0", x"56", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 3990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 367290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier =>       887,
         data => (x"25", x"51", x"75", x"15", x"b1", x"64", x"e0", x"80", x"74", x"40", x"b5", x"5d", x"ca", x"a6", x"c1", x"7f", x"97", x"1c", x"30", x"81", x"32", x"23", x"44", x"c0", x"63", x"9a", x"c6", x"35", x"9f", x"49", x"c7", x"44", x"1a", x"3e", x"d9", x"4c", x"a2", x"ba", x"4c", x"96", x"7b", x"02", x"74", x"46", x"28", x"36", x"45", x"bf", x"d1", x"f5", x"c1", x"04", x"19", x"06", x"44", x"7c", x"a0", x"0b", x"31", x"c0", x"d3", x"79", x"05", x"6e")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns),
           ('1', 251290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 305
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       975,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1690 ns), ('0', 2490 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 520810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       881,
         data => (x"db", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 516790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>       316,
         data => (x"17", x"32", x"71", x"af", x"b7", x"36", x"ab", x"59", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 339290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1575,
         data => (x"9e", x"04", x"0e", x"fd", x"3e", x"67", x"97", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 379290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1613,
         data => (x"88", x"fc", x"59", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 447290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1303,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1126,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 407817329,
         data => (x"d0", x"69", x"48", x"de", x"67", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 373310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1768,
         data => (x"ab", x"16", x"5c", x"34", x"14", x"35", x"5e", x"82", x"7b", x"1f", x"22", x"b3", x"0f", x"fa", x"21", x"ab", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 205310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 107
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>        24,
         data => (x"f5", x"e1", x"5d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 1490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 2010 ns),
           ('1', 504290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       439,
         data => (x"2d", x"3a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  28814705,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 10110 ns), ('0', 1990 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>        66,
         data => (x"7c", x"7a", x"34", x"f7", x"9c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 387310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 474868774,
         data => (x"03", x"fc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 10110 ns), ('0', 1990 ns), ('1', 423310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>  25430070,
         data => (x"eb", x"0f", x"f0", x"a5", x"04", x"b4", x"3c", x"ac", x"8c", x"08", x"33", x"e6", x"ce", x"58", x"e3", x"c9", x"8c", x"5b", x"66", x"6d", x"7f", x"53", x"f3", x"1c", x"d5", x"f0", x"1a", x"b6", x"c1", x"e1", x"7a", x"2e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 340310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 177
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 181407447,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       484,
         data => (x"15", x"e6", x"2b", x"78", x"b0", x"b8", x"d3", x"96", x"a5", x"53", x"e9", x"99", x"ef", x"c0", x"0a", x"89", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 207290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 97
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 258908507,
         data => (x"5c", x"5c", x"4e", x"50", x"fc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns),
           ('1', 460290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>   5407470,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 521030644,
         data => (x"a8", x"8b", x"24", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 403290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 492352006,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  52269070,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 478790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>      1208,
         data => (x"88", x"70", x"11", x"67", x"61", x"3c", x"5d", x"25", x"fb", x"3b", x"15", x"b3", x"c8", x"3d", x"3f", x"6d", x"8c", x"9d", x"fb", x"f4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 432790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 115
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 178640521,
         data => (x"27", x"88", x"c6", x"60", x"a8", x"d9", x"68", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 319310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1623,
         data => (x"2d", x"1f", x"a1", x"68", x"b4", x"55", x"b0", x"f1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 487790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>   1966107,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 474790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       203,
         data => (x"f3", x"81", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 435290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 459229266,
         data => (x"ca", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>  31926835,
         data => (x"c6", x"47", x"48", x"2f", x"fb", x"1e", x"60", x"6d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 293290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 198991537,
         data => (x"de", x"83", x"fb", x"39", x"e7", x"70", x"3a", x"d4", x"aa", x"9c", x"e9", x"bf", x"e6", x"98", x"40", x"80", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 163310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 109
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>  13216632,
         data => (x"f6", x"82", x"4c", x"d6", x"f0", x"fe", x"d5", x"dc", x"63", x"6d", x"3b", x"e7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 910 ns), ('0', 2010 ns), ('1', 430790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 91
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 428275352,
         data => (x"24", x"05", x"cb", x"8e", x"c4", x"b2", x"a6", x"84", x"b3", x"66", x"6a", x"7b", x"ed", x"99", x"72", x"70", x"65", x"c9", x"e0", x"e3", x"1f", x"bd", x"48", x"8c", x"79", x"30", x"75", x"6e", x"7f", x"4f", x"9d", x"24", x"d3", x"e9", x"b2", x"18", x"9c", x"59", x"9d", x"50", x"3f", x"87", x"cb", x"2d", x"a0", x"be", x"9e", x"86", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 2490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 2490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 281310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 239
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 140897602,
         data => (x"b2", x"33", x"37", x"62", x"a8", x"a5", x"62", x"77", x"c2", x"06", x"4b", x"ac", x"b8", x"64", x"c9", x"91", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 171310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 121
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1481,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1511,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>      1987,
         data => (x"4e", x"86", x"90", x"30", x"ae", x"b5", x"92", x"27", x"79", x"98", x"f1", x"a5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 468290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 91
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1746,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1540,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 185545236,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>  21548716,
         data => (x"1a", x"d4", x"56", x"48", x"0b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 460290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1581,
         data => (x"2a", x"d1", x"b7", x"1a", x"b4", x"10", x"24", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 383290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 168567778,
         data => (x"28", x"e6", x"38", x"68", x"d0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 345290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 498549374,
         data => (x"6a", x"8a", x"dd", x"75", x"72", x"cd", x"79", x"f3", x"2f", x"23", x"c6", x"e6", x"3d", x"fa", x"f6", x"e0", x"62", x"e7", x"f4", x"7b", x"e3", x"1d", x"62", x"9b", x"85", x"b2", x"2b", x"01", x"48", x"5f", x"96", x"32", x"e9", x"75", x"27", x"db", x"c2", x"20", x"d0", x"71", x"43", x"17", x"58", x"01", x"91", x"cf", x"e1", x"f3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 990 ns), ('0', 990 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 277310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 239
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       766,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       316,
         data => (x"7b", x"cb", x"42", x"13", x"7d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 500290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       780,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 1390 ns), ('0', 2010 ns), ('1', 520790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       697,
         data => (x"93", x"89", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 437290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 435417022,
         data => (x"42", x"63", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 391310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>       674,
         data => (x"b7", x"d2", x"ac", x"04", x"94", x"3f", x"81", x"c0", x"c6", x"a6", x"c8", x"90", x"6b", x"a1", x"4c", x"73", x"90", x"e0", x"fc", x"91", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 434310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 125
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 218918020,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       257,
         data => (x"12", x"54", x"d9", x"3f", x"d7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 2010 ns),
           ('1', 498290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1064,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 184732543,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>   7684517,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 453310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       904,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       118,
         data => (x"45", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 514810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 157982750,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1661,
         data => (x"cc", x"b3", x"bc", x"39", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 502810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1409,
         data => (x"f4", x"af", x"29", x"ba", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 433310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1351,
         data => (x"7a", x"5e", x"54", x"dd", x"f8", x"73", x"00", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 491790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1395,
         data => (x"07", x"84", x"6f", x"c3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 403310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1117,
         data => (x"85", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1085,
         data => (x"7f", x"30", x"e9", x"8e", x"2a", x"48", x"e3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 2010 ns),
           ('1', 492290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1917,
         data => (x"57", x"2a", x"e3", x"13", x"32", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 389290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>         0,
         data => (x"99", x"7c", x"70", x"9e", x"c7", x"d0", x"cd", x"cd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 335290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>        17,
         data => (x"a7", x"54", x"bf", x"30", x"15", x"96", x"b9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81900 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 383310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1038,
         data => (x"95", x"8d", x"05", x"0c", x"b3", x"c3", x"25", x"af", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1910 ns), ('0', 1990 ns),
           ('1', 486310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1523,
         data => (x"45", x"a6", x"5f", x"c2", x"b2", x"3b", x"ea", x"86", x"7b", x"1b", x"1b", x"91", x"d4", x"5c", x"00", x"39", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 205310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 97
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 142980578,
         data => (x"d9", x"42", x"c9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 470790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1743,
         data => (x"02", x"54", x"af", x"a9", x"33", x"f1", x"5c", x"6e", x"dc", x"63", x"69", x"78", x"7e", x"fb", x"4d", x"da", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 454310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 105
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       197,
         data => (x"ea", x"83", x"2e", x"ad", x"4d", x"ad", x"20", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 2010 ns),
           ('1', 491790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 263237046,
         data => (x"b9", x"f5", x"77", x"ac", x"d2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 349310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       851,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1147,
         data => (x"55", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 516810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1515,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       118,
         data => (x"5f", x"76", x"ae", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 506290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1842,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1326,
         data => (x"66", x"21", x"5e", x"31", x"70", x"6e", x"78", x"c5", x"da", x"3c", x"ef", x"32", x"04", x"c8", x"b6", x"98", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 211290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 99
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1618,
         data => (x"a3", x"00", x"f2", x"45", x"b1", x"88", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 399290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 366017389,
         data => (x"49", x"41", x"60", x"b9", x"30", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 375290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 271276569,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1423,
         data => (x"86", x"4f", x"aa", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 419290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1242,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 421133431,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 152260420,
         data => (x"56", x"7f", x"20", x"af", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 365310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 234533038,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       799,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>       534,
         data => (x"c4", x"50", x"1d", x"c2", x"a5", x"68", x"89", x"a3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 341310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>        24,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81900 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 495310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       247,
         data => (x"cb", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 483310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 386417810,
         data => (x"3e", x"28", x"bf", x"7c", x"21", x"43", x"86", x"65", x"13", x"24", x"28", x"b9", x"8c", x"b1", x"dc", x"24", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 416790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 111
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 211327790,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 459310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 528006817,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  79769664,
         data => (x"42", x"8f", x"b5", x"3e", x"b0", x"f9", x"45", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 335290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1335,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       632,
         data => (x"e8", x"45", x"a7", x"17", x"98", x"b3", x"2e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 355310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 318593955,
         data => (x"82", x"14", x"52", x"13", x"ca", x"10", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 333290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       186,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1651,
         data => (x"3a", x"4e", x"2a", x"a2", x"14", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 419290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       306,
         data => (x"e9", x"92", x"03", x"09", x"21", x"85", x"1d", x"73", x"18", x"e7", x"04", x"5c", x"2c", x"d8", x"b5", x"fd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 209290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 103
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1294,
         data => (x"4f", x"9a", x"02", x"f2", x"ae", x"54", x"2d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 491790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 255284656,
         data => (x"98", x"4e", x"8e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 409290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 419004385,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 451310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 204854098,
         data => (x"fc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 478310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 186590972,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 130050140,
         data => (x"c3", x"02", x"67", x"1f", x"17", x"ac", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 355290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 167127873,
         data => (x"e6", x"1c", x"03", x"3a", x"21", x"15", x"39", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 341310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 409155265,
         data => (x"49", x"38", x"e0", x"ab", x"96", x"51", x"01", x"23", x"94", x"82", x"0a", x"33", x"99", x"b7", x"3f", x"c8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 165290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 105
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 151377423,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 451290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 455614984,
         data => (x"15", x"8b", x"c4", x"8b", x"fe", x"8d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 357290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>      1739,
         data => (x"ba", x"fc", x"c5", x"3e", x"08", x"f8", x"57", x"bf", x"38", x"21", x"f1", x"11", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 263310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1604,
         data => (x"9a", x"fc", x"ec", x"b0", x"88", x"31", x"bb", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 383290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       870,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1445,
         data => (x"f1", x"de", x"d6", x"4a", x"1e", x"8e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 375310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 167565565,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 2010 ns), ('1', 427290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 174447012,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 8090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       697,
         data => (x"fd", x"d9", x"2c", x"65", x"d2", x"86", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 373290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       968,
         data => (x"bc", x"b0", x"c3", x"da", x"be", x"ae", x"6b", x"5f", x"cf", x"08", x"84", x"c0", x"05", x"44", x"ae", x"ee", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 205310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 99
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 183353035,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       518,
         data => (x"05", x"bd", x"70", x"de", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 431290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1144,
         data => (x"4e", x"2b", x"73", x"2d", x"fa", x"7b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 371290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier => 163820329,
         data => (x"ee", x"2b", x"8f", x"f8", x"8b", x"b1", x"db", x"19", x"3a", x"12", x"ab", x"3f", x"50", x"1c", x"9d", x"88", x"c8", x"2d", x"04", x"d0", x"fa", x"2f", x"44", x"29", x"aa", x"bf", x"5a", x"e5", x"41", x"50", x"50", x"30", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 345290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 195
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1873,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 189538579,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 459310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1712,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 379485725,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 371039414,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1824,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>      1948,
         data => (x"75", x"a5", x"46", x"c0", x"bc", x"92", x"cb", x"24", x"fa", x"73", x"14", x"ab", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 275290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 89
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 113862994,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 482790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 213043293,
         data => (x"2d", x"42", x"09", x"32", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 367310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  23866994,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 477058270,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier => 348858913,
         data => (x"77", x"cd", x"d3", x"7f", x"fb", x"ec", x"2b", x"f0", x"fe", x"a4", x"6b", x"e4", x"51", x"ae", x"6d", x"83", x"e8", x"95", x"99", x"44", x"e4", x"a3", x"45", x"79", x"ef", x"04", x"21", x"87", x"e7", x"43", x"14", x"de", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 346790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 187
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 244162553,
         data => (x"89", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 435310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       101,
         data => (x"fe", x"97", x"a6", x"83", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 427290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  77106008,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 467406759,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 9990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 453310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 189528921,
         data => (x"55", x"0f", x"34", x"b3", x"1c", x"89", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 335310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>         9,
         data => (x"96", x"6a", x"9b", x"3d", x"6d", x"1c", x"f8", x"89", x"61", x"9a", x"c9", x"6c", x"b4", x"f9", x"fa", x"70", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1990 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 453310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 103
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1083,
         data => (x"7c", x"b2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 435290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>      1014,
         data => (x"1a", x"23", x"36", x"30", x"8d", x"d1", x"6d", x"fa", x"6d", x"e5", x"04", x"ce", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 273290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 81
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>        13,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>       449,
         data => (x"79", x"ee", x"90", x"2d", x"e9", x"a8", x"e8", x"22", x"5b", x"82", x"45", x"91", x"b2", x"52", x"63", x"9f", x"cc", x"d0", x"86", x"d0", x"20", x"86", x"1e", x"da", x"3c", x"66", x"91", x"e1", x"61", x"39", x"f5", x"5b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 384790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 165
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1327,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 288463771,
         data => (x"1b", x"a6", x"cb", x"fd", x"c6", x"18", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 458290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>   1254428,
         data => (x"87", x"4a", x"90", x"6d", x"5c", x"f1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 357290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 479976298,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1814,
         data => (x"06", x"26", x"18", x"80", x"c1", x"3f", x"cb", x"bf", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1390 ns), ('0', 2010 ns), ('1', 486290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1518,
         data => (x"7d", x"26", x"d4", x"c8", x"36", x"43", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 397290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>      1317,
         data => (x"3d", x"78", x"fe", x"ef", x"c9", x"9b", x"93", x"4f", x"41", x"2c", x"cf", x"03", x"ea", x"1c", x"43", x"f0", x"01", x"d1", x"43", x"cd", x"50", x"69", x"a3", x"98", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 417810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 135
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1217,
         data => (x"76", x"d9", x"36", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 449310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 467729180,
         data => (x"39", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 437290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       954,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       356,
         data => (x"4f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 481310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       309,
         data => (x"b7", x"8d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 437310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 373173640,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 270479680,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 449290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  40286482,
         data => (x"bf", x"71", x"6e", x"0f", x"e4", x"ea", x"d0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 10010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 337290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 256160880,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       456,
         data => (x"04", x"25", x"14", x"ee", x"56", x"0f", x"48", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 351290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 100903158,
         data => (x"f2", x"14", x"48", x"64", x"02", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 371290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 263895677,
         data => (x"27", x"7c", x"3e", x"7f", x"3e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 367290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       686,
         data => (x"b2", x"22", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 211961364,
         data => (x"df", x"24", x"c7", x"69", x"17", x"5b", x"31", x"fa", x"dc", x"89", x"c3", x"4a", x"b1", x"66", x"71", x"ae", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 173310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 113
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       703,
         data => (x"f8", x"73", x"15", x"2b", x"16", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 498290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 304701218,
         data => (x"27", x"86", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 423310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1259,
         data => (x"18", x"1e", x"cb", x"db", x"68", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 419290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 102515362,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 480810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1793,
         data => (x"bf", x"df", x"bc", x"55", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 501790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier => 214320597,
         data => (x"c3", x"df", x"f2", x"d3", x"fc", x"34", x"15", x"15", x"d1", x"60", x"71", x"3a", x"5e", x"33", x"13", x"89", x"1a", x"5c", x"22", x"e5", x"27", x"b3", x"a6", x"07", x"ef", x"7b", x"fe", x"61", x"98", x"d7", x"70", x"db", x"b8", x"63", x"af", x"35", x"17", x"45", x"4b", x"e8", x"a5", x"3c", x"a2", x"83", x"ee", x"b5", x"0e", x"89", x"13", x"af", x"6f", x"3a", x"63", x"95", x"c1", x"53", x"12", x"40", x"35", x"2a", x"18", x"25", x"07", x"50")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1490 ns), ('0', 2490 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 216810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 319
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       926,
         data => (x"d1", x"88", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 465310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       416,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1463,
         data => (x"f5", x"ae", x"c5", x"8b", x"70", x"99", x"9d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 385290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 152297781,
         data => (x"cf", x"19", x"7b", x"85", x"9f", x"1b", x"02", x"f0", x"24", x"a3", x"7e", x"50", x"49", x"7a", x"31", x"fc", x"01", x"26", x"5f", x"f6", x"d4", x"26", x"82", x"c4", x"3f", x"21", x"f4", x"8d", x"69", x"bc", x"80", x"b8", x"d5", x"7b", x"3e", x"75", x"97", x"40", x"66", x"3b", x"e3", x"64", x"8b", x"ad", x"df", x"3c", x"2a", x"60", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 278290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 243
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 101939580,
         data => (x"59", x"fb", x"6e", x"f9", x"70", x"7b", x"63", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 311290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1529,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 347665406,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  39930494,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       360,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1198,
         data => (x"a8", x"fd", x"af", x"19", x"f9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 415290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1425,
         data => (x"6e", x"0a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 435310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 355817159,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 223896612,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1755,
         data => (x"ed", x"52", x"95", x"a3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 435310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       114,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 17
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1610,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 520810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1003,
         data => (x"12", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 514790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       456,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 8090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       710,
         data => (x"e1", x"8b", x"81", x"f6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       341,
         data => (x"97", x"e6", x"6e", x"9b", x"fb", x"96", x"0e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 353310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1697,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  25074908,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 364727145,
         data => (x"37", x"42", x"4a", x"ad", x"71", x"c7", x"b8", x"f2", x"d9", x"d0", x"5a", x"c7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 237290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 101
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 143713106,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       458,
         data => (x"0f", x"05", x"40", x"08", x"9f", x"59", x"5c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 7990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 377310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>  23150090,
         data => (x"c1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       669,
         data => (x"ca", x"58", x"d4", x"b7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 504790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 250892001,
         data => (x"2b", x"69", x"09", x"db", x"f7", x"0e", x"1c", x"7f", x"ae", x"75", x"5b", x"85", x"17", x"6f", x"9e", x"02", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 7990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 169310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 105
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>  13101048,
         data => (x"40", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 6110 ns), ('0', 2010 ns), ('1', 407290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1055,
         data => (x"48", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 512790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 141582715,
         data => (x"64", x"e5", x"2d", x"f2", x"03", x"2c", x"21", x"f7", x"87", x"a6", x"0f", x"76", x"45", x"91", x"27", x"ef", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 165290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 107
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       572,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 10110 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1772,
         data => (x"d4", x"94", x"3e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 508310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  32587588,
         data => (x"16", x"48", x"a2", x"37", x"c0", x"2b", x"dd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 311290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 167434571,
         data => (x"92", x"26", x"9b", x"aa", x"2d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 351290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 122683158,
         data => (x"ab", x"ae", x"22", x"e9", x"8e", x"6b", x"0d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 317290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>       494,
         data => (x"d9", x"5d", x"30", x"37", x"ad", x"52", x"da", x"0e", x"9b", x"ec", x"35", x"b6", x"98", x"e1", x"1b", x"dc", x"2a", x"f4", x"69", x"d5", x"a3", x"0b", x"3f", x"b2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 990 ns), ('0', 990 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 420310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 141
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 209943938,
         data => (x"24", x"de", x"4a", x"82", x"10", x"81", x"30", x"e1", x"5c", x"3e", x"fc", x"c9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 7990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 225310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 87
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 174747466,
         data => (x"be", x"7e", x"43", x"a7", x"d3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 373310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       850,
         data => (x"e0", x"20", x"83", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 198779456,
         data => (x"71", x"1d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 397310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier => 374677540,
         data => (x"c2", x"a8", x"03", x"a4", x"fc", x"51", x"e2", x"fb", x"14", x"0b", x"cf", x"7b", x"bd", x"63", x"14", x"67", x"c3", x"b4", x"6a", x"15", x"f9", x"4c", x"2f", x"41", x"3e", x"cb", x"38", x"91", x"c5", x"ec", x"e1", x"08", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 345790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 177
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       484,
         data => (x"8f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 525567469,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 453310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 331831634,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 2010 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 281090984,
         data => (x"4b", x"c9", x"34", x"17", x"02", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 349290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 311691956,
         data => (x"05", x"8c", x"92", x"18", x"43", x"22", x"27", x"0e", x"3d", x"85", x"d4", x"94", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 237290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 95
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 430539066,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 480790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1227,
         data => (x"11", x"26", x"cd", x"92", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 433310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 335533701,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 427290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier => 420824749,
         data => (x"c4", x"c4", x"71", x"02", x"ca", x"46", x"96", x"13", x"75", x"ea", x"62", x"b3", x"68", x"cd", x"fa", x"da", x"04", x"8b", x"81", x"51", x"1e", x"6d", x"7c", x"1f", x"00", x"0c", x"26", x"20", x"ae", x"c3", x"02", x"73", x"09", x"f2", x"f4", x"d3", x"b8", x"0b", x"66", x"ad", x"76", x"49", x"61", x"de", x"17", x"db", x"39", x"9a", x"67", x"ba", x"ec", x"85", x"28", x"e8", x"a5", x"29", x"74", x"4b", x"c8", x"a2", x"0f", x"ca", x"16", x"97")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 215810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 335
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier => 474759883,
         data => (x"d1", x"a5", x"0d", x"1b", x"86", x"6b", x"32", x"63", x"a4", x"4c", x"4a", x"60", x"39", x"50", x"88", x"a1", x"f5", x"31", x"17", x"c0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 990 ns), ('1', 990 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 990 ns), ('1', 910 ns), ('0', 2010 ns),
           ('1', 398290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 129
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       839,
         data => (x"e7", x"83", x"da", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 2510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1890 ns), ('0', 2010 ns),
           ('1', 507290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>      1836,
         data => (x"fd", x"3f", x"a6", x"69", x"f0", x"0a", x"8e", x"3e", x"d3", x"ee", x"f6", x"24", x"f6", x"19", x"99", x"29", x"30", x"5a", x"a2", x"69", x"aa", x"67", x"b9", x"92", x"ea", x"15", x"e4", x"e5", x"85", x"0a", x"05", x"04", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 385790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 175
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 410788223,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       851,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1593,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 329140052,
         data => (x"15", x"db", x"df", x"00", x"70", x"45", x"65", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 2010 ns),
           ('1', 311290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 409523680,
         data => (x"96", x"67", x"d1", x"cc", x"e3", x"c9", x"d6", x"cd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 301310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       669,
         data => (x"b9", x"f9", x"70", x"67", x"1c", x"bd", x"7c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 491310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 266223573,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 501329643,
         data => (x"c8", x"e3", x"41", x"1b", x"b0", x"a4", x"e4", x"07", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 301290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1259,
         data => (x"d8", x"5d", x"5a", x"49", x"c4", x"f5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 375290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1198,
         data => (x"d5", x"09", x"9e", x"b4", x"3a", x"eb", x"8e", x"03", x"d0", x"50", x"1e", x"01", x"f4", x"83", x"88", x"68", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 453790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 101
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 163415839,
         data => (x"e8", x"db", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 5990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 423310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1424,
         data => (x"bf", x"65", x"2a", x"95", x"ed", x"49", x"4b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 355310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1796,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 495310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>  88440930,
         data => (x"8f", x"07", x"ee", x"24", x"92", x"71", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 357290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 377746489,
         data => (x"1f", x"88", x"15", x"de", x"6d", x"40", x"f3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 337310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1308,
         data => (x"99", x"2f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 467290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  51176143,
         data => (x"46", x"da", x"e9", x"b4", x"fe", x"7c", x"a5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 317290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       226,
         data => (x"91", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 305698484,
         data => (x"64", x"2c", x"fe", x"24", x"30", x"bc", x"bd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 345290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1870,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 6110 ns), ('0', 2010 ns), ('1', 469290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       583,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 8090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      2019,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 6110 ns), ('0', 2010 ns),
           ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 17
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 189794320,
         data => (x"97", x"ec", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 391290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 495350134,
         data => (x"f4", x"a1", x"48", x"32", x"80", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 371290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>       483,
         data => (x"75", x"bd", x"e2", x"47", x"63", x"ab", x"bf", x"1a", x"6d", x"2a", x"2b", x"4f", x"a6", x"9f", x"66", x"13", x"e3", x"73", x"64", x"d4", x"fe", x"59", x"76", x"c6", x"0c", x"76", x"90", x"3f", x"ce", x"a7", x"55", x"44", x"65", x"38", x"8c", x"48", x"63", x"cb", x"63", x"d0", x"f6", x"8e", x"9f", x"1d", x"ad", x"06", x"31", x"92", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 321290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 239
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 191777354,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       949,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 493290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 455854551,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 474793690,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>  36179422,
         data => (x"1b", x"54", x"c4", x"a0", x"05", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 373290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      2024,
         data => (x"09", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 481290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 245280294,
         data => (x"bc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 441310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 304183305,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 254392895,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 234999219,
         data => (x"3d", x"fb", x"72", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 379290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1173,
         data => (x"1f", x"65", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 435310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       895,
         data => (x"a5", x"33", x"aa", x"ef", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 405290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier => 528116308,
         data => (x"bc", x"55", x"d9", x"f2", x"3e", x"12", x"c3", x"fa", x"0e", x"b5", x"bd", x"e1", x"42", x"1b", x"f2", x"e1", x"00", x"20", x"d2", x"e8", x"3f", x"e4", x"0e", x"72", x"0f", x"fe", x"23", x"2f", x"80", x"46", x"67", x"bd", x"1b", x"c1", x"b0", x"59", x"d3", x"f3", x"d4", x"61", x"aa", x"12", x"43", x"ec", x"ac", x"b5", x"ce", x"ad", x"d6", x"21", x"16", x"95", x"06", x"25", x"87", x"95", x"24", x"ab", x"c4", x"24", x"f1", x"ab", x"61", x"8d")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 2490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 2490 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 2490 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 210310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 305
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1678,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier =>       416,
         data => (x"1d", x"fa", x"1c", x"ec", x"28", x"72", x"8d", x"3f", x"08", x"14", x"64", x"8f", x"a9", x"08", x"3b", x"ed", x"2c", x"ad", x"19", x"0e", x"ba", x"07", x"9f", x"21", x"47", x"26", x"5d", x"e9", x"d6", x"2b", x"cf", x"f4", x"a5", x"eb", x"61", x"ce", x"5e", x"ee", x"0e", x"66", x"82", x"f1", x"75", x"2c", x"f9", x"31", x"1a", x"a5", x"5e", x"34", x"b3", x"19", x"ba", x"54", x"3a", x"02", x"f9", x"17", x"6c", x"51", x"c1", x"3c", x"46", x"68")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 252790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 303
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1560,
         data => (x"c4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 481290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       290,
         data => (x"30", x"12", x"df", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 447290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 379630972,
         data => (x"4e", x"dd", x"c3", x"50", x"d7", x"5a", x"3c", x"29", x"1d", x"78", x"ee", x"85", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 432810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 99
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  23773375,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 8110 ns), ('0', 2010 ns), ('1', 451290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       798,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 339974539,
         data => (x"76", x"7c", x"46", x"fe", x"ca", x"24", x"c2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 339290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 170713740,
         data => (x"ba", x"d0", x"95", x"bf", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 466310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 275412486,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 427290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       232,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  80931349,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 130455505,
         data => (x"42", x"d9", x"f2", x"be", x"f7", x"4b", x"65", x"32", x"1c", x"fa", x"f1", x"0c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 231290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 85
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 394650505,
         data => (x"cb", x"99", x"9d", x"e6", x"3f", x"38", x"88", x"4f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 303310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1851,
         data => (x"33", x"ef", x"90", x"27", x"ae", x"08", x"72", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 351310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 160217245,
         data => (x"1a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 8110 ns), ('0', 1990 ns), ('1', 441290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 495607931,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>        21,
         data => (x"d8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 479290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       408,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       788,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 168450362,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 8110 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       983,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 10090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 17
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1546,
         data => (x"72", x"8b", x"8b", x"62", x"97", x"e3", x"5b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 355290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier => 433706487,
         data => (x"44", x"15", x"65", x"25", x"27", x"18", x"0d", x"2a", x"df", x"30", x"bb", x"b6", x"fd", x"67", x"42", x"e5", x"50", x"81", x"d0", x"42", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 395310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 141
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  42411760,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 478790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 261879678,
         data => (x"6d", x"39", x"d5", x"52", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 460790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  37639569,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 8090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>       279,
         data => (x"c9", x"44", x"fe", x"99", x"c5", x"50", x"db", x"d1", x"2d", x"7f", x"75", x"ed", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 275290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 89
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       832,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 2010 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>  66082975,
         data => (x"a0", x"a6", x"f7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 405290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>      1740,
         data => (x"2d", x"f3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 463310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 162119019,
         data => (x"e8", x"ce", x"a8", x"68", x"44", x"97", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 337310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>       617,
         data => (x"7a", x"8a", x"c0", x"36", x"97", x"61", x"dc", x"8f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 488290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>        12,
         data => (x"50", x"c6", x"f9", x"fb", x"54", x"77", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 8110 ns), ('0', 2010 ns), ('1', 395290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 113412690,
         data => (x"0a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 439290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 190688628,
         data => (x"f7", x"46", x"76", x"b8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 393310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>       440,
         data => (x"43", x"28", x"bf", x"17", x"6a", x"10", x"dd", x"64", x"0d", x"b2", x"5b", x"85", x"6f", x"21", x"27", x"15", x"2b", x"60", x"23", x"05", x"2b", x"8e", x"fc", x"f0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 417810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 147
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 276587232,
         data => (x"47", x"ae", x"14", x"6f", x"6f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 5990 ns),
           ('1', 7990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 347290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1999,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 495310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 469063969,
         data => (x"3a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 413310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 314803656,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 9970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 229289169,
         data => (x"f6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 413310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>  33986921,
         data => (x"37", x"01", x"5a", x"26", x"ab", x"34", x"a5", x"b4", x"f1", x"31", x"f0", x"0b", x"43", x"1c", x"45", x"7c", x"5c", x"2a", x"95", x"40", x"14", x"d9", x"b2", x"fa", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 379290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 159
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       885,
         data => (x"83", x"1f", x"e9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 445310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1272,
         data => (x"35", x"e4", x"9e", x"67", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 500810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 208026879,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 5990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1169,
         data => (x"2d", x"95", x"41", x"a7", x"a6", x"6b", x"3f", x"d9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 487290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1133,
         data => (x"f2", x"97", x"77", x"a0", x"4c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 415310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       491,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       467,
         data => (x"f1", x"c0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 435310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1460,
         data => (x"fc", x"2b", x"86", x"d6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1371,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 536488145,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 349488222,
         data => (x"c6", x"b7", x"e4", x"4b", x"28", x"d6", x"8c", x"a6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 303290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 83
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 300371640,
         data => (x"91", x"42", x"b6", x"5a", x"0c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 2010 ns), ('1', 373290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>  16773439,
         data => (x"a4", x"30", x"45", x"89", x"d2", x"ad", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 450290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 71
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>   1450508,
         data => (x"3f", x"00", x"1b", x"4b", x"26", x"10", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 327310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 469869820,
         data => (x"0f", x"c5", x"f8", x"1b", x"cd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 369310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1965,
         data => (x"49", x"7a", x"66", x"1c", x"28", x"85", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 375290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1483,
         data => (x"dc", x"5a", x"27", x"03", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 405290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1083,
         data => (x"ae", x"46", x"2a", x"a7", x"e1", x"77", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 403290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       807,
         data => (x"5a", x"7b", x"5d", x"f6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       427,
         data => (x"32", x"9c", x"9c", x"0c", x"c4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 500290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       637,
         data => (x"7e", x"de", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 510290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>  92768331,
         data => (x"51", x"70", x"32", x"52", x"e6", x"0c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 455810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1116,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1870,
         data => (x"04", x"33", x"94", x"a3", x"aa", x"2f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 496310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       771,
         data => (x"56", x"b7", x"24", x"f7", x"0a", x"94", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 401290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 272778068,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81900 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 175020125,
         data => (x"50", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 194533962,
         data => (x"35", x"75", x"33", x"e3", x"c8", x"8c", x"11", x"7a", x"59", x"68", x"32", x"7e", x"df", x"bb", x"92", x"89", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 167290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 117
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       677,
         data => (x"78", x"df", x"35", x"27", x"30", x"03", x"7c", x"50", x"d4", x"85", x"05", x"c9", x"38", x"e8", x"12", x"44", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 453790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 103
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       742,
         data => (x"1d", x"c1", x"fa", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 417290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 258986458,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       628,
         data => (x"ab", x"66", x"c5", x"a7", x"36", x"1a", x"2d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 385290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>  47375006,
         data => (x"aa", x"9d", x"04", x"49", x"80", x"c2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 357310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 300234400,
         data => (x"52", x"54", x"19", x"a8", x"61", x"9c", x"de", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 452290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       553,
         data => (x"fa", x"83", x"9d", x"36", x"68", x"83", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 397290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       595,
         data => (x"f7", x"77", x"a4", x"5e", x"ba", x"63", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1910 ns), ('0', 1990 ns),
           ('1', 496790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1176,
         data => (x"dd", x"29", x"7d", x"bc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 2010 ns),
           ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1242,
         data => (x"fb", x"b8", x"d3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 508290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>      1868,
         data => (x"07", x"03", x"e1", x"7e", x"7b", x"06", x"dc", x"b5", x"69", x"50", x"7d", x"9e", x"18", x"5e", x"fb", x"41", x"5b", x"38", x"8d", x"a1", x"39", x"42", x"d7", x"35", x"fa", x"2c", x"e6", x"1b", x"84", x"72", x"1a", x"0b", x"f5", x"7b", x"89", x"f0", x"82", x"e6", x"a6", x"6b", x"37", x"a3", x"8a", x"50", x"02", x"86", x"11", x"5d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 317310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 237
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       228,
         data => (x"d6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 483290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 394285325,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  74924416,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 10110 ns), ('0', 1990 ns),
           ('1', 449290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1491,
         data => (x"94", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 516790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 244255744,
         data => (x"b9", x"8a", x"9b", x"96", x"c9", x"b9", x"95", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 315310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 73
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       477,
         data => (x"70", x"05", x"ec", x"78", x"8c", x"7d", x"0a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 2010 ns), ('1', 355290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 313060814,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>       945,
         data => (x"16", x"ec", x"fc", x"20", x"88", x"94", x"6a", x"c2", x"2a", x"2d", x"dd", x"97", x"9d", x"53", x"88", x"22", x"bf", x"80", x"af", x"bc", x"8a", x"39", x"c6", x"31", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 2490 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 418810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 133
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>  20392110,
         data => (x"bc", x"82", x"05", x"aa", x"7f", x"a4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 453310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1621,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 8090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1955,
         data => (x"dd", x"7c", x"66", x"5e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 504290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 270049919,
         data => (x"1b", x"17", x"48", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 405290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       163,
         data => (x"bb", x"dc", x"57", x"60", x"0f", x"eb", x"70", x"05", x"2a", x"2c", x"d7", x"7f", x"86", x"7e", x"5e", x"82", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 203290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 103
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       413,
         data => (x"13", x"f3", x"c0", x"aa", x"bb", x"b5", x"00", x"f2", x"e7", x"d7", x"2e", x"44", x"ae", x"8e", x"53", x"1a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 207310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 105
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>   9557767,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 478810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier => 483458122,
         data => (x"14", x"5e", x"62", x"9d", x"05", x"f4", x"11", x"45", x"9f", x"4c", x"fa", x"9f", x"be", x"62", x"f6", x"ec", x"a6", x"26", x"7c", x"7a", x"bf", x"fa", x"52", x"84", x"a6", x"03", x"48", x"58", x"32", x"6a", x"8c", x"46", x"48", x"6e", x"64", x"4d", x"64", x"f4", x"13", x"04", x"42", x"0e", x"24", x"01", x"71", x"1b", x"6e", x"97", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 2010 ns), ('1', 278290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 245
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1900,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 329534888,
         data => (x"e4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 478790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 379335641,
         data => (x"60", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 411290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1736,
         data => (x"49", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 451310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1616,
         data => (x"08", x"eb", x"f7", x"c9", x"56", x"89", x"ca", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 353290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 186566310,
         data => (x"1e", x"ac", x"70", x"d5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns),
           ('1', 385290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 188739642,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 453310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  17205564,
         data => (x"4c", x"f2", x"f9", x"c9", x"52", x"02", x"35", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 311290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 116488994,
         data => (x"c6", x"c2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 399310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1189,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 414926038,
         data => (x"58", x"f0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 399290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 105429886,
         data => (x"0d", x"48", x"a2", x"d7", x"1a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 375290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 143034337,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier =>      2024,
         data => (x"6c", x"15", x"ef", x"a7", x"1f", x"c9", x"80", x"79", x"78", x"58", x"6a", x"c9", x"f3", x"ab", x"9f", x"9c", x"b9", x"67", x"be", x"11", x"82", x"e3", x"1d", x"67", x"d3", x"35", x"20", x"59", x"93", x"1b", x"45", x"01", x"30", x"36", x"a8", x"4f", x"7f", x"a8", x"c9", x"f7", x"81", x"34", x"c1", x"75", x"60", x"e1", x"13", x"1a", x"49", x"d1", x"aa", x"cb", x"35", x"c7", x"b2", x"09", x"fd", x"52", x"e2", x"91", x"6e", x"28", x"12", x"1e")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 247790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 309
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1121,
         data => (x"37", x"55", x"65", x"ea", x"97", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 500810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 477442848,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 218998387,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       895,
         data => (x"e0", x"67", x"82", x"88", x"7a", x"a0", x"67", x"b4", x"0e", x"44", x"98", x"45", x"1a", x"7d", x"31", x"b1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 203290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 101
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>        87,
         data => (x"6d", x"84", x"71", x"7c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1741,
         data => (x"d2", x"d7", x"08", x"55", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 437290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 526083574,
         data => (x"84", x"0c", x"50", x"c9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 389290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       924,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 8110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1433,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 280849466,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       366,
         data => (x"bb", x"d2", x"98", x"bd", x"48", x"5f", x"75", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 1910 ns), ('0', 1990 ns), ('1', 492290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier => 477903709,
         data => (x"12", x"91", x"e8", x"b8", x"09", x"ea", x"a3", x"e1", x"5b", x"93", x"ac", x"c7", x"7d", x"41", x"72", x"5d", x"f4", x"ef", x"16", x"b1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 2470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 395290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 133
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 422625092,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       997,
         data => (x"8a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 479290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 443047592,
         data => (x"de", x"98", x"6b", x"3a", x"ab", x"97", x"81", x"a8", x"d8", x"f3", x"86", x"4e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 434290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 97
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 502513752,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 451290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       587,
         data => (x"d0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       407,
         data => (x"50", x"ad", x"80", x"ae", x"c5", x"6c", x"e9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 383310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier => 300528239,
         data => (x"df", x"a0", x"ab", x"c2", x"bc", x"2b", x"69", x"07", x"19", x"1a", x"de", x"6c", x"22", x"af", x"e9", x"19", x"8b", x"23", x"8f", x"5b", x"d1", x"90", x"0b", x"17", x"fc", x"74", x"09", x"80", x"5f", x"a4", x"5d", x"be", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1910 ns), ('0', 1990 ns),
           ('1', 347310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 185
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1400,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1105,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 520810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1606,
         data => (x"a3", x"47", x"cf", x"00", x"98", x"df", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 371290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 392103102,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 4110 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1673,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  34449694,
         data => (x"8a", x"ae", x"44", x"10", x"96", x"fd", x"b6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 9990 ns),
           ('1', 9990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 337310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1116,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 193281582,
         data => (x"30", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 413290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>  66897777,
         data => (x"c6", x"1c", x"56", x"e8", x"df", x"f5", x"0e", x"d6", x"80", x"bc", x"9b", x"10", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1910 ns), ('0', 1990 ns), ('1', 429810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 87
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1595,
         data => (x"3d", x"d4", x"23", x"04", x"a7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 500310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       337,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1464,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1052,
         data => (x"7a", x"62", x"67", x"b6", x"7d", x"f6", x"89", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 379290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1377,
         data => (x"df", x"f4", x"7f", x"87", x"18", x"2a", x"8b", x"eb", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 335310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>   1545146,
         data => (x"2b", x"14", x"f5", x"17", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 389290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 413765489,
         data => (x"c7", x"7f", x"ba", x"d0", x"16", x"78", x"dc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 343290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 295434445,
         data => (x"c4", x"75", x"9d", x"50", x"61", x"76", x"bc", x"88", x"5e", x"42", x"b3", x"72", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 432310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 97
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1706,
         data => (x"13", x"57", x"23", x"92", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 431290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 141931965,
         data => (x"11", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 441290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       691,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 138754079,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 5990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  61940457,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>       385,
         data => (x"a7", x"7b", x"c3", x"cb", x"8d", x"55", x"bf", x"b5", x"de", x"90", x"46", x"dc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 273310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 87
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 268068805,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 151021921,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 179304552,
         data => (x"ee", x"76", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 423290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>   8923406,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 339694363,
         data => (x"54", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 8090 ns), ('0', 2010 ns),
           ('1', 439290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       773,
         data => (x"fd", x"49", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 424794232,
         data => (x"d0", x"59", x"01", x"66", x"83", x"1c", x"d4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 7990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 313310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1188,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  17919659,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       679,
         data => (x"3e", x"31", x"49", x"08", x"85", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 2010 ns), ('1', 500290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1945,
         data => (x"0f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1705,
         data => (x"8c", x"9b", x"a3", x"25", x"ba", x"74", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 403290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 123799234,
         data => (x"d3", x"3a", x"45", x"1e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 393310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       744,
         data => (x"8a", x"66", x"b0", x"e9", x"1d", x"3f", x"c9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 383290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1440,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 220834626,
         data => (x"ac", x"81", x"7d", x"81", x"d2", x"51", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 331290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 157244298,
         data => (x"57", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 439290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier =>       597,
         data => (x"4c", x"b9", x"7b", x"96", x"f3", x"4d", x"5c", x"21", x"2c", x"bd", x"f0", x"b0", x"da", x"35", x"dd", x"5c", x"b3", x"de", x"af", x"84", x"9a", x"c7", x"74", x"50", x"56", x"4c", x"06", x"60", x"ae", x"a2", x"9c", x"7a", x"5d", x"97", x"90", x"51", x"e4", x"ec", x"f2", x"90", x"2b", x"e3", x"c1", x"06", x"99", x"9f", x"e1", x"cc", x"7e", x"91", x"d0", x"98", x"d8", x"46", x"68", x"af", x"92", x"ee", x"10", x"c0", x"91", x"ac", x"3b", x"6e")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 254290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 303
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier => 143067966,
         data => (x"33", x"b9", x"64", x"96", x"7b", x"e9", x"af", x"9a", x"cc", x"7c", x"98", x"dd", x"4e", x"31", x"b7", x"14", x"1a", x"67", x"26", x"09", x"77", x"e6", x"1a", x"a4", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 375290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 141
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1858,
         data => (x"11", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 516790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1200,
         data => (x"c5", x"76", x"c2", x"60", x"43", x"be", x"f8", x"a0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 2470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 485310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 67
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 339514717,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 237503188,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1959,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 5990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1422,
         data => (x"9e", x"f1", x"c7", x"64", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1910 ns), ('0', 2010 ns), ('1', 504790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 45
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  17507959,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 429290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       975,
         data => (x"f7", x"aa", x"63", x"3e", x"77", x"1a", x"6c", x"dd", x"75", x"bb", x"cd", x"39", x"f8", x"07", x"0d", x"de", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 209310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 101
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       614,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1071,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 495290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 440696597,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1415,
         data => (x"51", x"d0", x"f9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 419310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 503236608,
         data => (x"4e", x"0d", x"e3", x"0a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 359310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>        83,
         data => (x"9b", x"1f", x"cf", x"73", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 9990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 403290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>  25328180,
         data => (x"c7", x"cf", x"89", x"2c", x"6b", x"5b", x"fc", x"65", x"a2", x"88", x"ac", x"a2", x"8e", x"7a", x"af", x"f1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 2490 ns), ('0', 1490 ns), ('1', 2490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 412810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 113
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 300460813,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 459310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       467,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 499310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1232,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>      1717,
         data => (x"9b", x"b4", x"cc", x"3e", x"3d", x"f8", x"e0", x"4b", x"73", x"10", x"3e", x"77", x"f8", x"65", x"89", x"ab", x"f8", x"b6", x"fc", x"5d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 2470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 434290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 117
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       303,
         data => (x"f7", x"25", x"2a", x"b7", x"db", x"12", x"53", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 355290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 118828462,
         data => (x"71", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 415310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 270990288,
         data => (x"fa", x"3d", x"4c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns), ('1', 464290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 423167930,
         data => (x"5a", x"24", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 9970 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 4110 ns), ('0', 2010 ns),
           ('1', 423290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 456837147,
         data => (x"fa", x"05", x"f4", x"8d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 8110 ns), ('0', 2010 ns), ('1', 389290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1932,
         data => (x"c4", x"d9", x"6e", x"90", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 504790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       439,
         data => (x"a0", x"7d", x"3b", x"24", x"a1", x"50", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1890 ns), ('0', 2010 ns),
           ('1', 495790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>       771,
         data => (x"73", x"8b", x"12", x"f7", x"80", x"9f", x"cf", x"07", x"0c", x"b8", x"5b", x"50", x"92", x"ca", x"e1", x"ec", x"12", x"36", x"c3", x"16", x"56", x"c0", x"52", x"7a", x"62", x"22", x"78", x"a7", x"48", x"ea", x"bd", x"3b", x"76", x"cf", x"33", x"f7", x"ee", x"03", x"7e", x"fa", x"3b", x"da", x"cb", x"4d", x"a5", x"ad", x"3a", x"37", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 2510 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 319290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 241
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>      1274,
         data => (x"1f", x"b4", x"a0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 506310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 139636909,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>   4150466,
         data => (x"07", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 435310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>  69103171,
         data => (x"e0", x"8c", x"01", x"86", x"3a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 345310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1784,
         data => (x"d7", x"78", x"2a", x"0c", x"19", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 381310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       381,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       703,
         data => (x"68", x"05", x"28", x"6e", x"c6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 417290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>       740,
         data => (x"8d", x"99", x"92", x"aa", x"d3", x"9d", x"02", x"4c", x"47", x"0e", x"e4", x"b1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 277290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 87
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1703,
         data => (x"de", x"fa", x"6e", x"0e", x"64", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 2490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 499810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier => 103790087,
         data => (x"a2", x"0d", x"f1", x"f7", x"9a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 343290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       794,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 5990 ns), ('1', 4110 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 181814857,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       890,
         data => (x"86", x"a6", x"b2", x"74", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 435310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 481301258,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 429310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 331313133,
         data => (x"04", x"48", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 419290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 469119666,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>       392,
         data => (x"c7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 514790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier =>  75486873,
         data => (x"36", x"b1", x"68", x"ea", x"c7", x"cf", x"55", x"b1", x"70", x"d3", x"bd", x"1e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 235290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 99
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>      1699,
         data => (x"73", x"1b", x"89", x"47", x"a0", x"2f", x"f0", x"37", x"f6", x"b8", x"a4", x"86", x"b6", x"98", x"bc", x"e7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns),
           ('1', 454790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 105
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 316541538,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>  27418556,
         data => (x"16", x"e2", x"c6", x"d5", x"34", x"3a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 454790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 69
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 507495754,
         data => (x"f2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 10110 ns), ('0', 1990 ns), ('1', 437310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1599,
         data => (x"e1", x"05", x"28", x"4a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 502290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>        49,
         data => (x"5c", x"98", x"9e", x"7c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 403310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>  65367666,
         data => (x"14", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 439290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       787,
         data => (x"be", x"ec", x"53", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 508310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 461580689,
         data => (x"45", x"b7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 1990 ns),
           ('1', 395310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       426,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1829,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier =>       572,
         data => (x"0b", x"eb", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 433290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 505254860,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 27
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 259184468,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 359106978,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 186342115,
         data => (x"02", x"3b", x"59", x"98", x"6f", x"83", x"8f", x"e2", x"b7", x"1a", x"4e", x"65", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1890 ns), ('0', 2010 ns), ('1', 432790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 95
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1094,
         data => (x"2d", x"d1", x"f4", x"fa", x"20", x"5a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 4010 ns), ('1', 6090 ns), ('0', 2010 ns),
           ('1', 369290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>  52318148,
         data => (x"e9", x"6c", x"9a", x"eb", x"a8", x"f3", x"05", x"97", x"77", x"94", x"f9", x"ae", x"2f", x"48", x"94", x"26", x"fd", x"34", x"38", x"08", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 890 ns), ('0', 2010 ns), ('1', 393790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 131
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       593,
         data => (x"d6", x"69", x"50", x"59", x"55", x"86", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 890 ns), ('0', 2010 ns),
           ('1', 496290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 65
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1375,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1322,
         data => (x"dc", x"62", x"f0", x"2d", x"80", x"b3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 371310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 219888371,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1418,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 20, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1011", identifier =>       137,
         data => (x"46", x"f9", x"81", x"74", x"0f", x"a1", x"a3", x"b0", x"0c", x"cf", x"0d", x"6e", x"c0", x"3a", x"6f", x"74", x"eb", x"46", x"f2", x"82", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1910 ns), ('0', 2010 ns), ('1', 434790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 117
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>       907,
         data => (x"5d", x"d6", x"75", x"e0", x"d0", x"8b", x"27", x"4a", x"0d", x"1b", x"d8", x"2f", x"bf", x"89", x"3b", x"8f", x"16", x"29", x"cf", x"51", x"98", x"c3", x"bc", x"5f", x"36", x"3f", x"5c", x"6e", x"98", x"99", x"89", x"75", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 2490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 386810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 165
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>       513,
         data => (x"fd", x"8b", x"97", x"98", x"e3", x"c6", x"58", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 490290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier =>       428,
         data => (x"37", x"54", x"43", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 421310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  95460923,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>       919,
         data => (x"5e", x"89", x"a8", x"35", x"ca", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 417310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       853,
         data => (x"b9", x"92", x"a4", x"a6", x"93", x"0c", x"a9", x"3e", x"44", x"7e", x"82", x"3f", x"0f", x"a4", x"f0", x"df", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 7970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 205290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 101
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 483681189,
         data => (x"27", x"c5", x"62", x"db", x"90", x"16", x"0f", x"e5", x"e0", x"da", x"1f", x"f2", x"7f", x"c5", x"87", x"8b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns),
           ('1', 415310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 105
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  22124955,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>      1621,
         data => (x"90", x"10", x"a5", x"4d", x"4a", x"4c", x"92", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 10110 ns), ('0', 1990 ns), ('1', 387310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 333006659,
         data => (x"88", x"a3", x"92", x"a7", x"16", x"91", x"ec", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 910 ns), ('0', 2010 ns), ('1', 454790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 517460452,
         data => (x"c9", x"2b", x"7b", x"47", x"18", x"7b", x"a3", x"a8", x"8c", x"c8", x"75", x"56", x"15", x"08", x"03", x"bd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 173310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 119
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       468,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 6110 ns), ('0', 1990 ns), ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 440211607,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 183638191,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 431290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier => 204262112,
         data => (x"9c", x"d7", x"6d", x"a8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 367310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       630,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       930,
         data => (x"49", x"30", x"f1", x"a3", x"af", x"8c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 401290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 3, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0011", identifier => 350126870,
         data => (x"6a", x"fb", x"78", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 405290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       700,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1616,
         data => (x"5c", x"78", x"d2", x"cf", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 405310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 144511793,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 186222299,
         data => (x"c5", x"7d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 4090 ns), ('0', 2010 ns),
           ('1', 425290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier =>      1366,
         data => (x"f2", x"21", x"47", x"9a", x"a8", x"71", x"6b", x"cf", x"7e", x"bb", x"2c", x"f6", x"8e", x"fc", x"84", x"29", x"36", x"5c", x"f2", x"e1", x"d7", x"ec", x"9a", x"3e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns), ('1', 420290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 141
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 24, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1100", identifier => 250493958,
         data => (x"a4", x"cf", x"f1", x"45", x"96", x"0c", x"6d", x"08", x"78", x"3d", x"06", x"b3", x"69", x"fc", x"c2", x"e5", x"02", x"eb", x"1d", x"5e", x"5e", x"fe", x"b5", x"4b", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 376310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 147
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 431450412,
         data => (x"c2", x"30", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 4110 ns), ('0', 1990 ns),
           ('1', 397310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 344086586,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 4110 ns), ('0', 1990 ns), ('1', 455310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 201818246,
         data => (x"38", x"5a", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 468790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>      1836,
         data => (x"88", x"27", x"14", x"e7", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 2110 ns), ('0', 1990 ns),
           ('1', 433310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 41
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 207798859,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 459290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 48, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1110", identifier =>       250,
         data => (x"ad", x"86", x"c3", x"3d", x"af", x"72", x"3a", x"60", x"19", x"74", x"18", x"74", x"98", x"cd", x"91", x"22", x"83", x"9a", x"49", x"98", x"02", x"6e", x"e1", x"b4", x"ad", x"1f", x"e5", x"1f", x"02", x"5a", x"c0", x"30", x"e0", x"84", x"ec", x"90", x"77", x"28", x"f0", x"90", x"1c", x"0a", x"05", x"34", x"57", x"17", x"56", x"da", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1670 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns),
           ('1', 1970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns),
           ('1', 1470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1410 ns), ('0', 1990 ns), ('1', 317790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 235
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 12, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1001", identifier => 281306579,
         data => (x"55", x"67", x"bb", x"74", x"4e", x"da", x"f5", x"a8", x"9b", x"26", x"09", x"a0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 5990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 2490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 434310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 101
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>       619,
         data => (x"a8", x"57", x"14", x"ae", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 504790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 382574530,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 7990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  17111217,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>  70606694,
         data => (x"27", x"f8", x"87", x"c2", x"9e", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 9990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 8110 ns), ('0', 2010 ns), ('1', 369290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 47
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 4, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0100", identifier =>  99065423,
         data => (x"ed", x"b4", x"a4", x"c5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 393290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1020,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 497310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier =>  76840922,
         data => (x"38", x"c5", x"42", x"49", x"12", x"44", x"a9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1910 ns), ('0', 1990 ns), ('1', 452790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 175920289,
         data => (x"c1", x"5f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 4090 ns), ('0', 2010 ns), ('1', 421290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>  60866268,
         data => (x"7e", x"c2", x"68", x"51", x"94", x"9c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 357290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 57
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 179757850,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 5990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 7990 ns), ('1', 9990 ns), ('0', 3990 ns), ('1', 8110 ns), ('0', 1990 ns), ('1', 457310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>  66759727,
         data => (x"d5", x"50", x"23", x"0f", x"8d", x"d3", x"0b", x"e9", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 9970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 297290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 378972940,
         data => (x"76", x"20", x"c3", x"39", x"88", x"15", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 359290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier => 257909290,
         data => (x"76", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns),
           ('1', 476790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  23358877,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 8010 ns), ('1', 4090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       818,
         data => (x"ee", x"17", x"4a", x"58", x"2d", x"34", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 373290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       370,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 23
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 444461699,
         data => (x"7b", x"d0", x"e4", x"37", x"c6", x"f8", x"bc", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 9990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 5990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 7990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 9990 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 7990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns),
           ('1', 5990 ns), ('0', 5990 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 339310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       972,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier =>      1036,
         data => (x"0b", x"f5", x"16", x"3f", x"48", x"43", x"b7", x"10", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 9970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns),
           ('1', 1990 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 1990 ns), ('1', 6110 ns), ('0', 2010 ns), ('1', 335290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 63
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1498,
         data => (x"5f", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 453290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 39
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1365,
         data => (x"bd", x"57", x"4b", x"8f", x"24", x"d8", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 8010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 405290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 53
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 7, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0111", identifier => 459371997,
         data => (x"93", x"dd", x"66", x"29", x"9c", x"ae", x"6c", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 321290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 75
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1730,
         data => (x"e4", x"10", x"2f", x"48", x"a6", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 3990 ns),
           ('1', 2110 ns), ('0', 2010 ns), ('1', 415290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>      1045,
         data => (x"4e", x"c0", x"5e", x"a7", x"52", x"b1", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 6090 ns), ('0', 2010 ns), ('1', 371290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 61
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 257203586,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 6110 ns), ('0', 1990 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 8, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1000", identifier => 166226557,
         data => (x"f5", x"f4", x"76", x"bf", x"c3", x"5b", x"4f", x"f2", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 2470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 2010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 1410 ns), ('0', 1990 ns), ('1', 447290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 77
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 506674952,
         data => (x"17", x"c0", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 4010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 419290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 415667223,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 4110 ns), ('0', 1990 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 1, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0001", identifier =>      1176,
         data => (x"d3", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 10010 ns),
           ('1', 3970 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 910 ns), ('0', 2010 ns), ('1', 514790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 37
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 274491544,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 9990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 7990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 7990 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 2110 ns), ('0', 1990 ns), ('1', 427310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 43
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 361093524,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 10090 ns), ('0', 2010 ns), ('1', 457290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       406,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 21
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  91202705,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 33
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       514,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 2510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 910 ns), ('0', 1990 ns), ('1', 518790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 31
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '1', data_length => 64, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1111", identifier =>  89634545,
         data => (x"80", x"48", x"b8", x"75", x"f7", x"66", x"61", x"9d", x"0a", x"8b", x"86", x"89", x"85", x"e1", x"ad", x"f3", x"25", x"d7", x"5c", x"7e", x"c2", x"8b", x"af", x"cd", x"2a", x"0c", x"28", x"89", x"37", x"f5", x"8e", x"b7", x"bd", x"47", x"2e", x"b6", x"2d", x"0f", x"d3", x"b7", x"1a", x"d9", x"c0", x"9f", x"bb", x"6e", x"94", x"60", x"46", x"70", x"de", x"89", x"fc", x"8f", x"d6", x"27", x"1b", x"fe", x"31", x"52", x"75", x"bf", x"8a", x"33")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 1990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 7990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 2490 ns), ('1', 1490 ns), ('0', 1990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 990 ns), ('0', 2490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 1490 ns), ('0', 1990 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns),
           ('1', 2470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 1990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 990 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 990 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 970 ns), ('0', 510 ns), ('1', 1990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 490 ns),
           ('1', 1910 ns), ('0', 1990 ns), ('1', 214310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 323
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>       235,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 497290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 25
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier =>       170,
         data => (x"02", x"d2", x"9b", x"16", x"33", x"62", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 401290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 51
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier => 181540877,
         data => (x"42", x"2b", x"bc", x"41", x"db", x"8e", x"b6", x"9b", x"19", x"6a", x"a2", x"d1", x"53", x"d7", x"19", x"11", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 10010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 6010 ns),
           ('1', 1970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2090 ns), ('0', 2010 ns), ('1', 173290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 119
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>  52652811,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 7990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 6010 ns), ('1', 7990 ns), ('0', 1990 ns),
           ('1', 3990 ns), ('0', 1990 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 9990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 459310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 29
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '0', brs => '0', data_length => 6, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0110", identifier => 365353082,
         data => (x"19", x"c0", x"da", x"1d", x"e2", x"1d", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 6010 ns),
           ('1', 7970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns), ('1', 7970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 5970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 10010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 8010 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns), ('1', 1970 ns), ('0', 8010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 9970 ns), ('0', 8010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 3970 ns), ('0', 4010 ns), ('1', 2090 ns), ('0', 2010 ns),
           ('1', 359290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 49
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 5, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0101", identifier =>      1879,
         data => (x"15", x"be", x"c7", x"7f", x"62", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 5990 ns), ('0', 3990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1690 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 2490 ns), ('0', 990 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 1490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 1490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 990 ns), ('0', 990 ns),
           ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 910 ns), ('0', 1990 ns), ('1', 499810 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 59
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 16, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1010", identifier =>       972,
         data => (x"fc", x"ad", x"8a", x"6e", x"aa", x"84", x"7b", x"3d", x"32", x"6a", x"d5", x"72", x"45", x"72", x"d4", x"62", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 3990 ns), ('1', 7970 ns), ('0', 4010 ns), ('1', 3990 ns), ('0', 7990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1690 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 2490 ns), ('0', 490 ns),
           ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 990 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns), ('1', 490 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 1970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 490 ns), ('0', 990 ns), ('1', 490 ns), ('0', 1490 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 1490 ns), ('0', 990 ns), ('1', 470 ns), ('0', 510 ns), ('1', 990 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns), ('1', 990 ns), ('0', 990 ns), ('1', 1990 ns), ('0', 490 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns),
           ('1', 1910 ns), ('0', 1990 ns), ('1', 456310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 115
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '0', rtr => '0', brs => '1', data_length => 32, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "1101", identifier =>      1261,
         data => (x"d4", x"9c", x"6a", x"54", x"7e", x"83", x"27", x"38", x"36", x"0a", x"35", x"e3", x"94", x"a3", x"0e", x"99", x"1f", x"ca", x"4b", x"09", x"a1", x"3e", x"4e", x"93", x"13", x"30", x"4e", x"87", x"f0", x"2b", x"2a", x"c5", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 5970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1670 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 1010 ns), ('1', 1470 ns), ('0', 2510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1970 ns), ('0', 1510 ns), ('1', 1470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 1470 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 2470 ns), ('0', 510 ns),
           ('1', 970 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 2010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 2470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 2510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 2010 ns), ('1', 2470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 2510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1010 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 1510 ns),
           ('1', 470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 1510 ns), ('1', 970 ns), ('0', 1010 ns), ('1', 970 ns), ('0', 510 ns),
           ('1', 470 ns), ('0', 1510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1470 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns),
           ('1', 1470 ns), ('0', 510 ns), ('1', 970 ns), ('0', 510 ns), ('1', 470 ns), ('0', 510 ns), ('1', 1390 ns), ('0', 2010 ns),
           ('1', 385790 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 177
   ),
   (
    frame =>
        (frame_format => '1', ident_type => '1', rtr => '0', brs => '0', data_length => 2, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0010", identifier => 290506478,
         data => (x"41", x"fd", OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 5990 ns), ('1', 1990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 1990 ns),
           ('1', 1990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 3990 ns), ('1', 3990 ns), ('0', 5990 ns), ('1', 3990 ns), ('0', 1990 ns),
           ('1', 5970 ns), ('0', 2010 ns), ('1', 5990 ns), ('0', 3990 ns), ('1', 1970 ns), ('0', 10010 ns), ('1', 3970 ns), ('0', 4010 ns),
           ('1', 1990 ns), ('0', 9990 ns), ('1', 9990 ns), ('0', 1990 ns), ('1', 5990 ns), ('0', 1990 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 1990 ns), ('0', 3990 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns),
           ('1', 3970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 2110 ns), ('0', 1990 ns), ('1', 395310 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 55
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '0', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier =>      1456,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 2010 ns), ('1', 3970 ns), ('0', 8010 ns),
           ('1', 1970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 6010 ns),
           ('1', 6090 ns), ('0', 2010 ns), ('1', 499290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 19
   ),
   (
    frame =>
        (frame_format => '0', ident_type => '1', rtr => '1', brs => '0', data_length => 0, esi => '0', lbpf => '0',
         ivld => '0', lbtbi => 0, erf => '0', erf_pos => "0000", erf_erp => '0', erf_type => "000",
         timestamp => x"0000000000000000", rwcnt => 0, dlc => "0000", identifier => 183227647,
         data => (OTHERS => x"00")
        ),
    seq =>
        (
           ('1', 81920 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 5970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 2010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 1970 ns), ('0', 4010 ns), ('1', 9970 ns), ('0', 2010 ns), ('1', 7970 ns), ('0', 10010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 5970 ns), ('0', 4010 ns), ('1', 7970 ns), ('0', 2010 ns), ('1', 1970 ns), ('0', 4010 ns), ('1', 1970 ns), ('0', 2010 ns),
           ('1', 2090 ns), ('0', 2010 ns), ('1', 455290 ns),  OTHERS => ('1', 1 ns)
        ),
    seq_len => 35
   )
);
end package reference_data_set_5;

package body reference_data_set_5 is
end package body;
